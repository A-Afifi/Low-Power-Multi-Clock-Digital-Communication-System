module SYS_TOP (
	scan_clk, 
	scan_rst, 
	test_mode, 
	SE, 
	SI, 
	SO, 
	RST_N, 
	UART_CLK, 
	REF_CLK, 
	UART_RX_IN, 
	UART_TX_O, 
	parity_error, 
	framing_error);
   input scan_clk;
   input scan_rst;
   input test_mode;
   input SE;
   input [3:0] SI;
   output [3:0] SO;
   input RST_N;
   input UART_CLK;
   input REF_CLK;
   input UART_RX_IN;
   output UART_TX_O;
   output parity_error;
   output framing_error;

   // Internal wires
   wire FE_PHN10_n12__Exclude_0_NET;
   wire FE_PHN9_n10__Exclude_0_NET;
   wire FE_PHN8_n12__Exclude_0_NET;
   wire REF_CLK__L2_N0;
   wire REF_CLK__L1_N0;
   wire UART_CLK__L2_N0;
   wire UART_CLK__L1_N0;
   wire scan_clk__L12_N1;
   wire scan_clk__L12_N0;
   wire scan_clk__L11_N0;
   wire scan_clk__L10_N1;
   wire scan_clk__L10_N0;
   wire scan_clk__L9_N1;
   wire scan_clk__L9_N0;
   wire scan_clk__L8_N1;
   wire scan_clk__L8_N0;
   wire scan_clk__L7_N1;
   wire scan_clk__L7_N0;
   wire scan_clk__L6_N1;
   wire scan_clk__L6_N0;
   wire scan_clk__L5_N1;
   wire scan_clk__L5_N0;
   wire scan_clk__L4_N1;
   wire scan_clk__L4_N0;
   wire scan_clk__L3_N1;
   wire scan_clk__L3_N0;
   wire scan_clk__L2_N0;
   wire scan_clk__L1_N0;
   wire REF_CLK_M__L5_N15;
   wire REF_CLK_M__L5_N14;
   wire REF_CLK_M__L5_N13;
   wire REF_CLK_M__L5_N12;
   wire REF_CLK_M__L5_N11;
   wire REF_CLK_M__L5_N10;
   wire REF_CLK_M__L5_N9;
   wire REF_CLK_M__L5_N8;
   wire REF_CLK_M__L5_N7;
   wire REF_CLK_M__L5_N6;
   wire REF_CLK_M__L5_N5;
   wire REF_CLK_M__L5_N4;
   wire REF_CLK_M__L5_N3;
   wire REF_CLK_M__L5_N2;
   wire REF_CLK_M__L5_N1;
   wire REF_CLK_M__L5_N0;
   wire REF_CLK_M__L4_N3;
   wire REF_CLK_M__L4_N2;
   wire REF_CLK_M__L4_N1;
   wire REF_CLK_M__L4_N0;
   wire REF_CLK_M__L3_N1;
   wire REF_CLK_M__L3_N0;
   wire REF_CLK_M__L2_N0;
   wire REF_CLK_M__L1_N1;
   wire REF_CLK_M__L1_N0;
   wire Gated_ALU_CLK__L3_N0;
   wire Gated_ALU_CLK__L2_N0;
   wire Gated_ALU_CLK__L1_N0;
   wire UART_CLK_M__L13_N0;
   wire UART_CLK_M__L12_N0;
   wire UART_CLK_M__L11_N0;
   wire UART_CLK_M__L10_N0;
   wire UART_CLK_M__L9_N0;
   wire UART_CLK_M__L8_N0;
   wire UART_CLK_M__L7_N1;
   wire UART_CLK_M__L7_N0;
   wire UART_CLK_M__L6_N1;
   wire UART_CLK_M__L6_N0;
   wire UART_CLK_M__L5_N1;
   wire UART_CLK_M__L5_N0;
   wire UART_CLK_M__L4_N0;
   wire UART_CLK_M__L3_N0;
   wire UART_CLK_M__L2_N1;
   wire UART_CLK_M__L2_N0;
   wire UART_CLK_M__L1_N0;
   wire n10__Exclude_0_NET;
   wire n12__Exclude_0_NET;
   wire RX_CLK_M__L3_N1;
   wire RX_CLK_M__L3_N0;
   wire RX_CLK_M__L2_N0;
   wire RX_CLK_M__L1_N0;
   wire TX_CLK_M__L3_N3;
   wire TX_CLK_M__L3_N2;
   wire TX_CLK_M__L3_N1;
   wire TX_CLK_M__L3_N0;
   wire TX_CLK_M__L2_N0;
   wire TX_CLK_M__L1_N0;
   wire FE_OFN7_SE;
   wire FE_OFN5_M_Domain2_SYNC_RST;
   wire FE_OFN4_M_Domain1_SYNC_RST;
   wire FE_OFN2_M_Domain1_SYNC_RST;
   wire FE_OFN1_M_Domain1_SYNC_RST;
   wire FE_OFN0_M_Domain1_SYNC_RST;
   wire REF_CLK_M;
   wire UART_CLK_M;
   wire RX_CLK;
   wire RX_CLK_M;
   wire TX_CLK;
   wire TX_CLK_M;
   wire M_RST_N;
   wire Domain1_SYNC_RST;
   wire M_Domain1_SYNC_RST;
   wire Domain2_SYNC_RST;
   wire M_Domain2_SYNC_RST;
   wire Sync_Valid;
   wire Rd_D_Valid_RF;
   wire RdEn_RF;
   wire WrEn_RF;
   wire ALU_OUT_Valid;
   wire ALU_EN;
   wire FIFO_FULL;
   wire WR_INC;
   wire CLK_Gating_EN;
   wire RX_OUT_Valid;
   wire TX_Busy;
   wire TX_IN_Valid;
   wire RD_INC;
   wire _1_net_;
   wire Gated_ALU_CLK;
   wire n2;
   wire n3;
   wire n4;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n17;
   wire n19;
   wire n20;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire [7:0] Sync_Data;
   wire [7:0] Rd_D_RF;
   wire [3:0] Addr_RF;
   wire [7:0] Wr_D_RF;
   wire [15:0] ALU_OUT;
   wire [3:0] ALU_FUN;
   wire [7:0] WR_Data;
   wire [7:0] DIV_RATIO;
   wire [3:0] RX_Div_Ratio;
   wire [7:0] UART_Config;
   wire [7:0] RX_OUT;
   wire [7:0] TX_IN;
   wire [7:0] Op_A;
   wire [7:0] Op_B;

   assign SO[2] = ALU_OUT[7] ;

   BUFX2M FE_PHC10_n12__Exclude_0_NET (.Y(FE_PHN8_n12__Exclude_0_NET), 
	.A(FE_PHN10_n12__Exclude_0_NET));
   DLY4X1M FE_PHC9_n10__Exclude_0_NET (.Y(n10__Exclude_0_NET), 
	.A(FE_PHN9_n10__Exclude_0_NET));
   DLY3X1M FE_PHC8_n12__Exclude_0_NET (.Y(n12__Exclude_0_NET), 
	.A(FE_PHN8_n12__Exclude_0_NET));
   CLKINVX40M REF_CLK__L2_I0 (.Y(REF_CLK__L2_N0), 
	.A(REF_CLK__L1_N0));
   CLKINVX40M REF_CLK__L1_I0 (.Y(REF_CLK__L1_N0), 
	.A(REF_CLK));
   CLKINVX40M UART_CLK__L2_I0 (.Y(UART_CLK__L2_N0), 
	.A(UART_CLK__L1_N0));
   CLKINVX40M UART_CLK__L1_I0 (.Y(UART_CLK__L1_N0), 
	.A(UART_CLK));
   CLKBUFX12M scan_clk__L12_I1 (.Y(scan_clk__L12_N1), 
	.A(scan_clk__L11_N0));
   CLKBUFX24M scan_clk__L12_I0 (.Y(scan_clk__L12_N0), 
	.A(scan_clk__L11_N0));
   CLKBUFX24M scan_clk__L11_I0 (.Y(scan_clk__L11_N0), 
	.A(scan_clk__L10_N1));
   CLKBUFX24M scan_clk__L10_I1 (.Y(scan_clk__L10_N1), 
	.A(scan_clk__L9_N1));
   BUFX8M scan_clk__L10_I0 (.Y(scan_clk__L10_N0), 
	.A(scan_clk__L9_N0));
   CLKBUFX24M scan_clk__L9_I1 (.Y(scan_clk__L9_N1), 
	.A(scan_clk__L8_N1));
   CLKBUFX24M scan_clk__L9_I0 (.Y(scan_clk__L9_N0), 
	.A(scan_clk__L8_N0));
   CLKBUFX24M scan_clk__L8_I1 (.Y(scan_clk__L8_N1), 
	.A(scan_clk__L7_N1));
   CLKBUFX24M scan_clk__L8_I0 (.Y(scan_clk__L8_N0), 
	.A(scan_clk__L7_N0));
   CLKBUFX24M scan_clk__L7_I1 (.Y(scan_clk__L7_N1), 
	.A(scan_clk__L6_N1));
   CLKBUFX24M scan_clk__L7_I0 (.Y(scan_clk__L7_N0), 
	.A(scan_clk__L6_N0));
   CLKBUFX24M scan_clk__L6_I1 (.Y(scan_clk__L6_N1), 
	.A(scan_clk__L5_N1));
   CLKBUFX24M scan_clk__L6_I0 (.Y(scan_clk__L6_N0), 
	.A(scan_clk__L5_N0));
   CLKBUFX24M scan_clk__L5_I1 (.Y(scan_clk__L5_N1), 
	.A(scan_clk__L4_N1));
   CLKBUFX24M scan_clk__L5_I0 (.Y(scan_clk__L5_N0), 
	.A(scan_clk__L4_N0));
   CLKBUFX24M scan_clk__L4_I1 (.Y(scan_clk__L4_N1), 
	.A(scan_clk__L3_N1));
   CLKBUFX24M scan_clk__L4_I0 (.Y(scan_clk__L4_N0), 
	.A(scan_clk__L3_N0));
   BUFX8M scan_clk__L3_I1 (.Y(scan_clk__L3_N1), 
	.A(scan_clk__L2_N0));
   BUFX12M scan_clk__L3_I0 (.Y(scan_clk__L3_N0), 
	.A(scan_clk__L2_N0));
   CLKINVX24M scan_clk__L2_I0 (.Y(scan_clk__L2_N0), 
	.A(scan_clk__L1_N0));
   CLKINVX40M scan_clk__L1_I0 (.Y(scan_clk__L1_N0), 
	.A(scan_clk));
   CLKINVX40M REF_CLK_M__L5_I15 (.Y(REF_CLK_M__L5_N15), 
	.A(REF_CLK_M__L4_N3));
   CLKINVX40M REF_CLK_M__L5_I14 (.Y(REF_CLK_M__L5_N14), 
	.A(REF_CLK_M__L4_N3));
   CLKINVX40M REF_CLK_M__L5_I13 (.Y(REF_CLK_M__L5_N13), 
	.A(REF_CLK_M__L4_N3));
   CLKINVX40M REF_CLK_M__L5_I12 (.Y(REF_CLK_M__L5_N12), 
	.A(REF_CLK_M__L4_N3));
   CLKINVX40M REF_CLK_M__L5_I11 (.Y(REF_CLK_M__L5_N11), 
	.A(REF_CLK_M__L4_N2));
   CLKINVX40M REF_CLK_M__L5_I10 (.Y(REF_CLK_M__L5_N10), 
	.A(REF_CLK_M__L4_N2));
   CLKINVX40M REF_CLK_M__L5_I9 (.Y(REF_CLK_M__L5_N9), 
	.A(REF_CLK_M__L4_N2));
   CLKINVX40M REF_CLK_M__L5_I8 (.Y(REF_CLK_M__L5_N8), 
	.A(REF_CLK_M__L4_N2));
   CLKINVX40M REF_CLK_M__L5_I7 (.Y(REF_CLK_M__L5_N7), 
	.A(REF_CLK_M__L4_N1));
   CLKINVX40M REF_CLK_M__L5_I6 (.Y(REF_CLK_M__L5_N6), 
	.A(REF_CLK_M__L4_N1));
   CLKINVX40M REF_CLK_M__L5_I5 (.Y(REF_CLK_M__L5_N5), 
	.A(REF_CLK_M__L4_N1));
   CLKINVX40M REF_CLK_M__L5_I4 (.Y(REF_CLK_M__L5_N4), 
	.A(REF_CLK_M__L4_N1));
   CLKINVX40M REF_CLK_M__L5_I3 (.Y(REF_CLK_M__L5_N3), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX40M REF_CLK_M__L5_I2 (.Y(REF_CLK_M__L5_N2), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX40M REF_CLK_M__L5_I1 (.Y(REF_CLK_M__L5_N1), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX40M REF_CLK_M__L5_I0 (.Y(REF_CLK_M__L5_N0), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX40M REF_CLK_M__L4_I3 (.Y(REF_CLK_M__L4_N3), 
	.A(REF_CLK_M__L3_N1));
   CLKINVX40M REF_CLK_M__L4_I2 (.Y(REF_CLK_M__L4_N2), 
	.A(REF_CLK_M__L3_N1));
   CLKINVX40M REF_CLK_M__L4_I1 (.Y(REF_CLK_M__L4_N1), 
	.A(REF_CLK_M__L3_N0));
   CLKINVX40M REF_CLK_M__L4_I0 (.Y(REF_CLK_M__L4_N0), 
	.A(REF_CLK_M__L3_N0));
   CLKINVX40M REF_CLK_M__L3_I1 (.Y(REF_CLK_M__L3_N1), 
	.A(REF_CLK_M__L2_N0));
   CLKINVX40M REF_CLK_M__L3_I0 (.Y(REF_CLK_M__L3_N0), 
	.A(REF_CLK_M__L2_N0));
   CLKINVX40M REF_CLK_M__L2_I0 (.Y(REF_CLK_M__L2_N0), 
	.A(REF_CLK_M__L1_N0));
   BUFX32M REF_CLK_M__L1_I1 (.Y(REF_CLK_M__L1_N1), 
	.A(REF_CLK_M));
   CLKBUFX12M REF_CLK_M__L1_I0 (.Y(REF_CLK_M__L1_N0), 
	.A(REF_CLK_M));
   CLKINVX32M Gated_ALU_CLK__L3_I0 (.Y(Gated_ALU_CLK__L3_N0), 
	.A(Gated_ALU_CLK__L2_N0));
   BUFX14M Gated_ALU_CLK__L2_I0 (.Y(Gated_ALU_CLK__L2_N0), 
	.A(Gated_ALU_CLK__L1_N0));
   CLKINVX6M Gated_ALU_CLK__L1_I0 (.Y(Gated_ALU_CLK__L1_N0), 
	.A(Gated_ALU_CLK));
   CLKINVX40M UART_CLK_M__L13_I0 (.Y(UART_CLK_M__L13_N0), 
	.A(UART_CLK_M__L12_N0));
   CLKINVX40M UART_CLK_M__L12_I0 (.Y(UART_CLK_M__L12_N0), 
	.A(UART_CLK_M__L11_N0));
   CLKBUFX40M UART_CLK_M__L11_I0 (.Y(UART_CLK_M__L11_N0), 
	.A(UART_CLK_M__L10_N0));
   CLKBUFX24M UART_CLK_M__L10_I0 (.Y(UART_CLK_M__L10_N0), 
	.A(UART_CLK_M__L9_N0));
   CLKBUFX24M UART_CLK_M__L9_I0 (.Y(UART_CLK_M__L9_N0), 
	.A(UART_CLK_M__L8_N0));
   CLKBUFX24M UART_CLK_M__L8_I0 (.Y(UART_CLK_M__L8_N0), 
	.A(UART_CLK_M__L7_N1));
   CLKBUFX24M UART_CLK_M__L7_I1 (.Y(UART_CLK_M__L7_N1), 
	.A(UART_CLK_M__L6_N1));
   CLKBUFX24M UART_CLK_M__L7_I0 (.Y(UART_CLK_M__L7_N0), 
	.A(UART_CLK_M__L6_N0));
   CLKBUFX24M UART_CLK_M__L6_I1 (.Y(UART_CLK_M__L6_N1), 
	.A(UART_CLK_M__L5_N1));
   CLKBUFX24M UART_CLK_M__L6_I0 (.Y(UART_CLK_M__L6_N0), 
	.A(UART_CLK_M__L5_N0));
   CLKBUFX24M UART_CLK_M__L5_I1 (.Y(UART_CLK_M__L5_N1), 
	.A(UART_CLK_M__L4_N0));
   BUFX14M UART_CLK_M__L5_I0 (.Y(UART_CLK_M__L5_N0), 
	.A(UART_CLK_M__L4_N0));
   CLKBUFX24M UART_CLK_M__L4_I0 (.Y(UART_CLK_M__L4_N0), 
	.A(UART_CLK_M__L3_N0));
   CLKBUFX24M UART_CLK_M__L3_I0 (.Y(UART_CLK_M__L3_N0), 
	.A(UART_CLK_M__L2_N0));
   BUFX8M UART_CLK_M__L2_I1 (.Y(UART_CLK_M__L2_N1), 
	.A(UART_CLK_M__L1_N0));
   CLKBUFX24M UART_CLK_M__L2_I0 (.Y(UART_CLK_M__L2_N0), 
	.A(UART_CLK_M__L1_N0));
   CLKBUFX12M UART_CLK_M__L1_I0 (.Y(UART_CLK_M__L1_N0), 
	.A(UART_CLK_M));
   BUFX8M n10__Exclude_0 (.Y(FE_PHN9_n10__Exclude_0_NET), 
	.A(n10));
   BUFX8M n12__Exclude_0 (.Y(FE_PHN10_n12__Exclude_0_NET), 
	.A(n12));
   CLKINVX32M RX_CLK_M__L3_I1 (.Y(RX_CLK_M__L3_N1), 
	.A(RX_CLK_M__L2_N0));
   CLKINVX32M RX_CLK_M__L3_I0 (.Y(RX_CLK_M__L3_N0), 
	.A(RX_CLK_M__L2_N0));
   CLKINVX32M RX_CLK_M__L2_I0 (.Y(RX_CLK_M__L2_N0), 
	.A(RX_CLK_M__L1_N0));
   CLKBUFX12M RX_CLK_M__L1_I0 (.Y(RX_CLK_M__L1_N0), 
	.A(RX_CLK_M));
   CLKINVX24M TX_CLK_M__L3_I3 (.Y(TX_CLK_M__L3_N3), 
	.A(TX_CLK_M__L2_N0));
   CLKINVX24M TX_CLK_M__L3_I2 (.Y(TX_CLK_M__L3_N2), 
	.A(TX_CLK_M__L2_N0));
   CLKINVX24M TX_CLK_M__L3_I1 (.Y(TX_CLK_M__L3_N1), 
	.A(TX_CLK_M__L2_N0));
   CLKINVX24M TX_CLK_M__L3_I0 (.Y(TX_CLK_M__L3_N0), 
	.A(TX_CLK_M__L2_N0));
   CLKINVX40M TX_CLK_M__L2_I0 (.Y(TX_CLK_M__L2_N0), 
	.A(TX_CLK_M__L1_N0));
   CLKBUFX20M TX_CLK_M__L1_I0 (.Y(TX_CLK_M__L1_N0), 
	.A(TX_CLK_M));
   BUFX4M FE_OFC7_SE (.Y(FE_OFN7_SE), 
	.A(SE));
   BUFX5M FE_OFC5_M_Domain2_SYNC_RST (.Y(FE_OFN5_M_Domain2_SYNC_RST), 
	.A(M_Domain2_SYNC_RST));
   CLKINVX6M FE_OFC4_M_Domain1_SYNC_RST (.Y(FE_OFN4_M_Domain1_SYNC_RST), 
	.A(FE_OFN0_M_Domain1_SYNC_RST));
   CLKINVX8M FE_OFC2_M_Domain1_SYNC_RST (.Y(FE_OFN2_M_Domain1_SYNC_RST), 
	.A(FE_OFN0_M_Domain1_SYNC_RST));
   CLKINVX6M FE_OFC1_M_Domain1_SYNC_RST (.Y(FE_OFN1_M_Domain1_SYNC_RST), 
	.A(FE_OFN0_M_Domain1_SYNC_RST));
   CLKINVX1M FE_OFC0_M_Domain1_SYNC_RST (.Y(FE_OFN0_M_Domain1_SYNC_RST), 
	.A(M_Domain1_SYNC_RST));
   OR2X2M U5 (.Y(_1_net_), 
	.B(n2), 
	.A(CLK_Gating_EN));
   BUFX2M U6 (.Y(n3), 
	.A(Addr_RF[0]));
   BUFX4M U7 (.Y(n4), 
	.A(Addr_RF[1]));
   BUFX2M U11 (.Y(n2), 
	.A(test_mode));
   DLY1X4M U14 (.Y(n25), 
	.A(n26));
   INVXLM U15 (.Y(n26), 
	.A(n34));
   DLY1X4M U16 (.Y(n27), 
	.A(n29));
   INVXLM U17 (.Y(n28), 
	.A(n37));
   INVXLM U18 (.Y(n29), 
	.A(n28));
   DLY1X4M U19 (.Y(n30), 
	.A(n37));
   DLY1X1M U20 (.Y(n31), 
	.A(n37));
   INVXLM U21 (.Y(n32), 
	.A(n36));
   CLKINVX2M U22 (.Y(n33), 
	.A(n32));
   INVXLM U23 (.Y(n34), 
	.A(FE_OFN7_SE));
   CLKINVX2M U24 (.Y(n35), 
	.A(n34));
   INVXLM U25 (.Y(n36), 
	.A(n34));
   CLKINVX2M U26 (.Y(n37), 
	.A(n34));
   mux2X1_1 DFT_REF_MUX (.IN_0(REF_CLK__L2_N0), 
	.IN_1(scan_clk__L10_N0), 
	.SEL(n2), 
	.OUT(REF_CLK_M));
   mux2X1_4 UART_CLK_MUX (.IN_0(UART_CLK__L2_N0), 
	.IN_1(scan_clk__L2_N0), 
	.SEL(n2), 
	.OUT(UART_CLK_M));
   mux2X1_3 RX_CLK_MUX (.IN_0(RX_CLK), 
	.IN_1(scan_clk__L12_N1), 
	.SEL(n2), 
	.OUT(RX_CLK_M));
   mux2X1_2 TX_CLK_MUX (.IN_0(TX_CLK), 
	.IN_1(scan_clk__L12_N0), 
	.SEL(n2), 
	.OUT(TX_CLK_M));
   mux2X1_0 RST_N_MUX (.IN_0(RST_N), 
	.IN_1(scan_rst), 
	.SEL(n2), 
	.OUT(M_RST_N));
   mux2X1_6 Domain1_SYNC_RST_MUX (.IN_0(Domain1_SYNC_RST), 
	.IN_1(scan_rst), 
	.SEL(n2), 
	.OUT(M_Domain1_SYNC_RST));
   mux2X1_5 Domain2_SYNC_RST_MUX (.IN_0(Domain2_SYNC_RST), 
	.IN_1(scan_rst), 
	.SEL(n2), 
	.OUT(M_Domain2_SYNC_RST));
   SYS_CTRL_D_Width8_Addr_Size4_test_1 SYS_Cntroller (.CLK(REF_CLK_M__L5_N1), 
	.RST(M_Domain1_SYNC_RST), 
	.Sync_Frame({ Sync_Data[7],
		Sync_Data[6],
		Sync_Data[5],
		Sync_Data[4],
		Sync_Data[3],
		Sync_Data[2],
		Sync_Data[1],
		Sync_Data[0] }), 
	.enable_pulse(Sync_Valid), 
	.Rd_D({ Rd_D_RF[7],
		Rd_D_RF[6],
		Rd_D_RF[5],
		Rd_D_RF[4],
		Rd_D_RF[3],
		Rd_D_RF[2],
		Rd_D_RF[1],
		Rd_D_RF[0] }), 
	.Rd_D_Valid(Rd_D_Valid_RF), 
	.Rd_En(RdEn_RF), 
	.Wr_En(WrEn_RF), 
	.Addr({ Addr_RF[3],
		Addr_RF[2],
		Addr_RF[1],
		Addr_RF[0] }), 
	.Wr_D({ Wr_D_RF[7],
		Wr_D_RF[6],
		Wr_D_RF[5],
		Wr_D_RF[4],
		Wr_D_RF[3],
		Wr_D_RF[2],
		Wr_D_RF[1],
		Wr_D_RF[0] }), 
	.ALU_OUT({ ALU_OUT[15],
		ALU_OUT[14],
		ALU_OUT[13],
		ALU_OUT[12],
		ALU_OUT[11],
		ALU_OUT[10],
		ALU_OUT[9],
		ALU_OUT[8],
		ALU_OUT[7],
		ALU_OUT[6],
		ALU_OUT[5],
		ALU_OUT[4],
		ALU_OUT[3],
		ALU_OUT[2],
		ALU_OUT[1],
		ALU_OUT[0] }), 
	.OUT_Valid(ALU_OUT_Valid), 
	.ALU_En(ALU_EN), 
	.FUN({ ALU_FUN[3],
		ALU_FUN[2],
		ALU_FUN[1],
		ALU_FUN[0] }), 
	.FIFO_FULL(FIFO_FULL), 
	.WR_INC(WR_INC), 
	.WR_DATA({ WR_Data[7],
		WR_Data[6],
		WR_Data[5],
		WR_Data[4],
		WR_Data[3],
		WR_Data[2],
		WR_Data[1],
		WR_Data[0] }), 
	.Gate_En(CLK_Gating_EN), 
	.test_si(n20), 
	.test_so(n19), 
	.test_se(n27), 
	.FE_OFN1_M_Domain1_SYNC_RST(FE_OFN1_M_Domain1_SYNC_RST), 
	.FE_OFN2_M_Domain1_SYNC_RST(FE_OFN2_M_Domain1_SYNC_RST), 
	.FE_OFN4_M_Domain1_SYNC_RST(FE_OFN4_M_Domain1_SYNC_RST), 
	.REF_CLK_M__L5_N14(REF_CLK_M__L5_N14), 
	.REF_CLK_M__L5_N2(REF_CLK_M__L5_N2), 
	.REF_CLK_M__L5_N3(REF_CLK_M__L5_N3));
   Integer_ClkDiv_ratio_Width8_test_1 UART_TX_ClkDiv (.i_ref_clk(UART_CLK_M__L13_N0), 
	.i_rst_n(M_Domain2_SYNC_RST), 
	.i_clk_en(1'b1), 
	.i_div_ratio({ DIV_RATIO[7],
		DIV_RATIO[6],
		DIV_RATIO[5],
		DIV_RATIO[4],
		DIV_RATIO[3],
		DIV_RATIO[2],
		DIV_RATIO[1],
		DIV_RATIO[0] }), 
	.o_div_clk(TX_CLK), 
	.test_si(n11), 
	.test_so(n10), 
	.test_se(n37), 
	.UART_CLK_M__L1_N0(UART_CLK_M__L1_N0), 
	.UART_CLK_M__L6_N1(UART_CLK_M__L6_N1));
   Integer_ClkDiv_ratio_Width4_test_1 UART_RX_ClkDiv (.i_ref_clk(UART_CLK_M__L13_N0), 
	.i_rst_n(FE_OFN5_M_Domain2_SYNC_RST), 
	.i_clk_en(1'b1), 
	.i_div_ratio({ RX_Div_Ratio[3],
		RX_Div_Ratio[2],
		RX_Div_Ratio[1],
		RX_Div_Ratio[0] }), 
	.o_div_clk(RX_CLK), 
	.test_si(n13), 
	.test_so(n12), 
	.test_se(n37), 
	.UART_CLK_M__L2_N1(UART_CLK_M__L2_N1), 
	.UART_CLK_M__L7_N0(UART_CLK_M__L7_N0));
   RX_CLKDIV_MUX_Width4 CLKDIV_MUX (.Input({ UART_Config[7],
		UART_Config[6],
		UART_Config[5],
		UART_Config[4],
		UART_Config[3],
		UART_Config[2] }), 
	.MUX_Out({ RX_Div_Ratio[3],
		RX_Div_Ratio[2],
		RX_Div_Ratio[1],
		RX_Div_Ratio[0] }));
   UART_RX_TOP_Data_Width8_test_1 UART_RX (.CLK(RX_CLK_M__L3_N0), 
	.RST(M_Domain2_SYNC_RST), 
	.PAR_EN(UART_Config[0]), 
	.Prescale({ UART_Config[7],
		UART_Config[6],
		UART_Config[5],
		UART_Config[4],
		UART_Config[3],
		UART_Config[2] }), 
	.PAR_TYP(UART_Config[1]), 
	.RX_IN(UART_RX_IN), 
	.Paerity_Error(parity_error), 
	.Stop_Error(framing_error), 
	.Data_Valid(RX_OUT_Valid), 
	.P_DATA({ RX_OUT[7],
		RX_OUT[6],
		RX_OUT[5],
		RX_OUT[4],
		RX_OUT[3],
		RX_OUT[2],
		RX_OUT[1],
		RX_OUT[0] }), 
	.test_si(Domain2_SYNC_RST), 
	.test_so(n13), 
	.test_se(n25), 
	.FE_OFN5_M_Domain2_SYNC_RST(FE_OFN5_M_Domain2_SYNC_RST), 
	.RX_CLK_M__L3_N1(RX_CLK_M__L3_N1));
   UART_TOP_test_1 UART_TX (.CLK(TX_CLK_M__L3_N0), 
	.RST(M_Domain2_SYNC_RST), 
	.P_DATA({ TX_IN[7],
		TX_IN[6],
		TX_IN[5],
		TX_IN[4],
		TX_IN[3],
		TX_IN[2],
		TX_IN[1],
		TX_IN[0] }), 
	.Data_Valid(TX_IN_Valid), 
	.PAR_EN(UART_Config[0]), 
	.PAR_TYP(UART_Config[1]), 
	.busy(TX_Busy), 
	.TX_OUT(SO[0]), 
	.test_si2(n10__Exclude_0_NET), 
	.test_si1(n12__Exclude_0_NET), 
	.test_so1(n11), 
	.test_se(n30), 
	.FE_OFN5_M_Domain2_SYNC_RST(FE_OFN5_M_Domain2_SYNC_RST), 
	.TX_CLK_M__L3_N1(TX_CLK_M__L3_N1), 
	.TX_CLK_M__L3_N2(TX_CLK_M__L3_N2), 
	.TX_CLK_M__L3_N3(TX_CLK_M__L3_N3));
   AS_FIFO_TOP_Data_Width8_Addr_Size3_FIFO_Dipth8_NUM_STAGES2_test_1 UART_FIFO (.I_W_CLK(REF_CLK_M__L5_N0), 
	.I_W_RST(M_Domain1_SYNC_RST), 
	.I_W_INC(WR_INC), 
	.I_Data({ WR_Data[7],
		WR_Data[6],
		WR_Data[5],
		WR_Data[4],
		WR_Data[3],
		WR_Data[2],
		WR_Data[1],
		WR_Data[0] }), 
	.I_R_CLK(TX_CLK_M__L3_N2), 
	.I_R_RST(M_Domain2_SYNC_RST), 
	.I_R_INC(RD_INC), 
	.O_Data({ TX_IN[7],
		TX_IN[6],
		TX_IN[5],
		TX_IN[4],
		TX_IN[3],
		TX_IN[2],
		TX_IN[1],
		TX_IN[0] }), 
	.FIFO_Full(FIFO_FULL), 
	.FIFO_Empty(TX_IN_Valid), 
	.test_si2(SI[0]), 
	.test_si1(n17), 
	.test_so2(n14), 
	.test_so1(SO[1]), 
	.test_se(FE_OFN7_SE), 
	.FE_OFN1_M_Domain1_SYNC_RST(FE_OFN1_M_Domain1_SYNC_RST), 
	.FE_OFN4_M_Domain1_SYNC_RST(FE_OFN4_M_Domain1_SYNC_RST), 
	.FE_OFN5_M_Domain2_SYNC_RST(FE_OFN5_M_Domain2_SYNC_RST), 
	.TX_CLK_M__L3_N3(TX_CLK_M__L3_N3), 
	.REF_CLK_M__L5_N1(REF_CLK_M__L5_N1), 
	.REF_CLK_M__L5_N4(REF_CLK_M__L5_N4), 
	.REF_CLK_M__L5_N5(REF_CLK_M__L5_N5), 
	.REF_CLK_M__L5_N6(REF_CLK_M__L5_N6), 
	.REF_CLK_M__L5_N7(REF_CLK_M__L5_N7));
   PULSE_GEN_test_1 U0_PULSE_GEN (.clk(TX_CLK_M__L3_N0), 
	.rst(M_Domain2_SYNC_RST), 
	.lvl_sig(TX_Busy), 
	.pulse_sig(RD_INC), 
	.test_si(ALU_OUT_Valid), 
	.test_so(n17), 
	.test_se(n31));
   RST_SYN_NUM_STAGES2_test_0 REF_RST_SYNC (.RST(M_RST_N), 
	.CLK(REF_CLK_M__L5_N0), 
	.SYNC_RST(Domain1_SYNC_RST), 
	.test_si(Sync_Data[7]), 
	.test_se(n33));
   RST_SYN_NUM_STAGES2_test_1 UART_RST_SYNC (.RST(M_RST_N), 
	.CLK(UART_CLK_M__L13_N0), 
	.SYNC_RST(Domain2_SYNC_RST), 
	.test_si(n14), 
	.test_se(n33));
   DATA_SYNC_NUM_STAGES2_BUS_WIDTH8_test_1 Data_SYNC (.CLK(REF_CLK_M__L5_N0), 
	.RST(M_Domain1_SYNC_RST), 
	.unsync_bus({ RX_OUT[7],
		RX_OUT[6],
		RX_OUT[5],
		RX_OUT[4],
		RX_OUT[3],
		RX_OUT[2],
		RX_OUT[1],
		RX_OUT[0] }), 
	.bus_enable(RX_OUT_Valid), 
	.sync_bus({ Sync_Data[7],
		Sync_Data[6],
		Sync_Data[5],
		Sync_Data[4],
		Sync_Data[3],
		Sync_Data[2],
		Sync_Data[1],
		Sync_Data[0] }), 
	.enable_pulse_d(Sync_Valid), 
	.test_si(SI[3]), 
	.test_se(n33), 
	.REF_CLK_M__L5_N2(REF_CLK_M__L5_N2), 
	.REF_CLK_M__L5_N3(REF_CLK_M__L5_N3));
   CLK_GATE U_CLK_GATE (.CLK_EN(_1_net_), 
	.CLK(REF_CLK_M__L1_N1), 
	.GATED_CLK(Gated_ALU_CLK));
   ALU_IN_Width8_test_1 U0_ALU (.CLK(Gated_ALU_CLK__L3_N0), 
	.RST(FE_OFN1_M_Domain1_SYNC_RST), 
	.EN(ALU_EN), 
	.ALU_FUN({ ALU_FUN[3],
		ALU_FUN[2],
		ALU_FUN[1],
		ALU_FUN[0] }), 
	.A({ Op_A[7],
		Op_A[6],
		Op_A[5],
		Op_A[4],
		Op_A[3],
		Op_A[2],
		Op_A[1],
		Op_A[0] }), 
	.B({ Op_B[7],
		Op_B[6],
		Op_B[5],
		Op_B[4],
		Op_B[3],
		Op_B[2],
		Op_B[1],
		Op_B[0] }), 
	.ALU_OUT({ ALU_OUT[15],
		ALU_OUT[14],
		ALU_OUT[13],
		ALU_OUT[12],
		ALU_OUT[11],
		ALU_OUT[10],
		ALU_OUT[9],
		ALU_OUT[8],
		ALU_OUT[7],
		ALU_OUT[6],
		ALU_OUT[5],
		ALU_OUT[4],
		ALU_OUT[3],
		ALU_OUT[2],
		ALU_OUT[1],
		ALU_OUT[0] }), 
	.OUT_Valid(ALU_OUT_Valid), 
	.test_si2(SI[1]), 
	.test_si1(n19), 
	.test_se(n35), 
	.FE_OFN4_M_Domain1_SYNC_RST(FE_OFN4_M_Domain1_SYNC_RST));
   Reg_File_WIDTH8_DEPTH16_ADDR4_test_1 RegFile (.CLK(REF_CLK_M__L5_N10), 
	.RST(FE_OFN0_M_Domain1_SYNC_RST), 
	.WrEn(WrEn_RF), 
	.RdEn(RdEn_RF), 
	.Address({ Addr_RF[3],
		Addr_RF[2],
		n4,
		n3 }), 
	.WrData({ Wr_D_RF[7],
		Wr_D_RF[6],
		Wr_D_RF[5],
		Wr_D_RF[4],
		Wr_D_RF[3],
		Wr_D_RF[2],
		Wr_D_RF[1],
		Wr_D_RF[0] }), 
	.RdData({ Rd_D_RF[7],
		Rd_D_RF[6],
		Rd_D_RF[5],
		Rd_D_RF[4],
		Rd_D_RF[3],
		Rd_D_RF[2],
		Rd_D_RF[1],
		Rd_D_RF[0] }), 
	.RdData_VLD(Rd_D_Valid_RF), 
	.REG0({ Op_A[7],
		Op_A[6],
		Op_A[5],
		Op_A[4],
		Op_A[3],
		Op_A[2],
		Op_A[1],
		Op_A[0] }), 
	.REG1({ Op_B[7],
		Op_B[6],
		Op_B[5],
		Op_B[4],
		Op_B[3],
		Op_B[2],
		Op_B[1],
		Op_B[0] }), 
	.REG2({ UART_Config[7],
		UART_Config[6],
		UART_Config[5],
		UART_Config[4],
		UART_Config[3],
		UART_Config[2],
		UART_Config[1],
		UART_Config[0] }), 
	.REG3({ DIV_RATIO[7],
		DIV_RATIO[6],
		DIV_RATIO[5],
		DIV_RATIO[4],
		DIV_RATIO[3],
		DIV_RATIO[2],
		DIV_RATIO[1],
		DIV_RATIO[0] }), 
	.test_si2(SI[2]), 
	.test_si1(Domain1_SYNC_RST), 
	.test_so2(n20), 
	.test_so1(SO[3]), 
	.test_se(FE_OFN7_SE), 
	.FE_OFN2_M_Domain1_SYNC_RST(FE_OFN2_M_Domain1_SYNC_RST), 
	.FE_OFN4_M_Domain1_SYNC_RST(FE_OFN4_M_Domain1_SYNC_RST), 
	.REF_CLK_M__L5_N11(REF_CLK_M__L5_N11), 
	.REF_CLK_M__L5_N12(REF_CLK_M__L5_N12), 
	.REF_CLK_M__L5_N13(REF_CLK_M__L5_N13), 
	.REF_CLK_M__L5_N14(REF_CLK_M__L5_N14), 
	.REF_CLK_M__L5_N15(REF_CLK_M__L5_N15), 
	.REF_CLK_M__L5_N3(REF_CLK_M__L5_N3), 
	.REF_CLK_M__L5_N8(REF_CLK_M__L5_N8), 
	.REF_CLK_M__L5_N9(REF_CLK_M__L5_N9));
   BUFX2M U13 (.Y(UART_TX_O), 
	.A(SO[0]));
endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : K-2015.06
// Date      : Wed Oct  1 07:11:59 2025
/////////////////////////////////////////////////////////////
module mux2X1_1 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   MX2X6M U1 (.Y(OUT), 
	.S0(N0), 
	.B(IN_1), 
	.A(IN_0));
endmodule

module mux2X1_4 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   MX2X2M U1 (.Y(OUT), 
	.S0(N0), 
	.B(IN_1), 
	.A(IN_0));
endmodule

module mux2X1_3 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   MX2X2M U1 (.Y(OUT), 
	.S0(N0), 
	.B(IN_1), 
	.A(IN_0));
endmodule

module mux2X1_2 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   MX2X2M U1 (.Y(OUT), 
	.S0(N0), 
	.B(IN_1), 
	.A(IN_0));
endmodule

module mux2X1_0 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   // Internal wires
   wire FE_PHN5_scan_rst;
   wire FE_PHN2_scan_rst;
   wire FE_PHN1_RST_N;
   wire FE_PHN0_RST_N;
   wire N0;

   assign N0 = SEL ;

   DLY4X1M FE_PHC5_scan_rst (.Y(FE_PHN5_scan_rst), 
	.A(FE_PHN2_scan_rst));
   DLY4X1M FE_PHC2_scan_rst (.Y(FE_PHN2_scan_rst), 
	.A(IN_1));
   DLY4X1M FE_PHC1_RST_N (.Y(FE_PHN1_RST_N), 
	.A(FE_PHN0_RST_N));
   DLY4X1M FE_PHC0_RST_N (.Y(FE_PHN0_RST_N), 
	.A(IN_0));
   MX2X2M U1 (.Y(OUT), 
	.S0(N0), 
	.B(FE_PHN5_scan_rst), 
	.A(FE_PHN1_RST_N));
endmodule

module mux2X1_6 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   // Internal wires
   wire FE_PHN6_scan_rst;
   wire FE_PHN3_scan_rst;
   wire N0;

   assign N0 = SEL ;

   DLY4X1M FE_PHC6_scan_rst (.Y(FE_PHN6_scan_rst), 
	.A(FE_PHN3_scan_rst));
   DLY4X1M FE_PHC3_scan_rst (.Y(FE_PHN3_scan_rst), 
	.A(IN_1));
   MX2X6M U1 (.Y(OUT), 
	.S0(N0), 
	.B(FE_PHN6_scan_rst), 
	.A(IN_0));
endmodule

module mux2X1_5 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   // Internal wires
   wire FE_PHN7_scan_rst;
   wire FE_PHN4_scan_rst;
   wire N0;

   assign N0 = SEL ;

   DLY4X1M FE_PHC7_scan_rst (.Y(FE_PHN7_scan_rst), 
	.A(FE_PHN4_scan_rst));
   DLY4X1M FE_PHC4_scan_rst (.Y(FE_PHN4_scan_rst), 
	.A(IN_1));
   CLKMX2X6M U1 (.Y(OUT), 
	.S0(N0), 
	.B(FE_PHN7_scan_rst), 
	.A(IN_0));
endmodule

module SYS_CTRL_D_Width8_Addr_Size4_test_1 (
	CLK, 
	RST, 
	Sync_Frame, 
	enable_pulse, 
	Rd_D, 
	Rd_D_Valid, 
	Rd_En, 
	Wr_En, 
	Addr, 
	Wr_D, 
	ALU_OUT, 
	OUT_Valid, 
	ALU_En, 
	FUN, 
	FIFO_FULL, 
	WR_INC, 
	WR_DATA, 
	Gate_En, 
	CLK_DIV_EN, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN1_M_Domain1_SYNC_RST, 
	FE_OFN2_M_Domain1_SYNC_RST, 
	FE_OFN4_M_Domain1_SYNC_RST, 
	REF_CLK_M__L5_N14, 
	REF_CLK_M__L5_N2, 
	REF_CLK_M__L5_N3);
   input CLK;
   input RST;
   input [7:0] Sync_Frame;
   input enable_pulse;
   input [7:0] Rd_D;
   input Rd_D_Valid;
   output Rd_En;
   output Wr_En;
   output [3:0] Addr;
   output [7:0] Wr_D;
   input [15:0] ALU_OUT;
   input OUT_Valid;
   output ALU_En;
   output [3:0] FUN;
   input FIFO_FULL;
   output WR_INC;
   output [7:0] WR_DATA;
   output Gate_En;
   output CLK_DIV_EN;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN1_M_Domain1_SYNC_RST;
   input FE_OFN2_M_Domain1_SYNC_RST;
   input FE_OFN4_M_Domain1_SYNC_RST;
   input REF_CLK_M__L5_N14;
   input REF_CLK_M__L5_N2;
   input REF_CLK_M__L5_N3;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n50;
   wire n54;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n48;
   wire n49;
   wire n51;
   wire n52;
   wire n53;
   wire n55;
   wire n56;
   wire n57;
   wire n66;
   wire n67;
   wire n68;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire [3:0] current_state;
   wire [3:0] next_state;
   wire [7:0] Stored_Frame1;

   assign test_so = current_state[3] ;

   TIELOM LTIE_LTIELO (.Y(LTIE_LTIELO_NET));
   SDFFRX1M \Stored_Frame2_reg[7]  (.SI(n160), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n40), 
	.Q(n159), 
	.D(n137), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRX1M \Stored_Frame2_reg[6]  (.SI(n161), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n41), 
	.Q(n160), 
	.D(n138), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRX1M \Stored_Frame2_reg[5]  (.SI(n162), 
	.SE(test_se), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.QN(n42), 
	.Q(n161), 
	.D(n139), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRX1M \Stored_Frame2_reg[4]  (.SI(n163), 
	.SE(test_se), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.QN(n43), 
	.Q(n162), 
	.D(n140), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRX1M \Stored_Frame3_reg[7]  (.SI(n152), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n58), 
	.Q(n151), 
	.D(n129), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRX1M \Stored_Frame3_reg[6]  (.SI(n153), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n59), 
	.Q(n152), 
	.D(n128), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRX1M \Stored_Frame3_reg[5]  (.SI(n154), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n60), 
	.Q(n153), 
	.D(n127), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRX1M \Stored_Frame3_reg[4]  (.SI(n155), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n61), 
	.Q(n154), 
	.D(n126), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRX1M \Stored_Frame3_reg[3]  (.SI(n156), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n62), 
	.Q(n155), 
	.D(n125), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRX1M \Stored_Frame3_reg[2]  (.SI(n157), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n63), 
	.Q(n156), 
	.D(n124), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRX1M \Stored_Frame3_reg[1]  (.SI(n158), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n64), 
	.Q(n157), 
	.D(n123), 
	.CK(CLK));
   SDFFRX1M \Stored_Frame3_reg[0]  (.SI(n159), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n65), 
	.Q(n158), 
	.D(n122), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRX1M \Stored_Frame1_reg[3]  (.SI(n148), 
	.SE(test_se), 
	.RN(RST), 
	.QN(n54), 
	.Q(n168), 
	.D(n134), 
	.CK(CLK));
   SDFFRQX2M \Stored_Frame1_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(Stored_Frame1[0]), 
	.D(n145), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \Stored_Frame1_reg[4]  (.SI(n168), 
	.SE(test_se), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(Stored_Frame1[4]), 
	.D(n133), 
	.CK(CLK));
   SDFFRX1M \Stored_Frame2_reg[3]  (.SI(n164), 
	.SE(test_se), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.QN(n44), 
	.Q(n163), 
	.D(n141), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRX1M \Stored_Frame2_reg[2]  (.SI(n165), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n45), 
	.Q(n164), 
	.D(n142), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRX1M \Stored_Frame2_reg[1]  (.SI(n166), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n46), 
	.Q(n165), 
	.D(n143), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \current_state_reg[0]  (.SI(n151), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(current_state[0]), 
	.D(next_state[0]), 
	.CK(CLK));
   SDFFRQX2M \Stored_Frame1_reg[6]  (.SI(Stored_Frame1[5]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Stored_Frame1[6]), 
	.D(n131), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \Stored_Frame1_reg[5]  (.SI(n147), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Stored_Frame1[5]), 
	.D(n132), 
	.CK(CLK));
   SDFFRQX2M \Stored_Frame1_reg[2]  (.SI(Stored_Frame1[1]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Stored_Frame1[2]), 
	.D(n135), 
	.CK(CLK));
   SDFFRQX2M \Stored_Frame1_reg[1]  (.SI(n57), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Stored_Frame1[1]), 
	.D(n136), 
	.CK(CLK));
   SDFFRX1M \Stored_Frame2_reg[0]  (.SI(n167), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n47), 
	.Q(n166), 
	.D(n144), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \current_state_reg[1]  (.SI(n150), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(current_state[1]), 
	.D(next_state[1]), 
	.CK(CLK));
   SDFFRQX2M \current_state_reg[3]  (.SI(n73), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(current_state[3]), 
	.D(next_state[3]), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \current_state_reg[2]  (.SI(n72), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(current_state[2]), 
	.D(next_state[2]), 
	.CK(CLK));
   SDFFRX1M \Stored_Frame1_reg[7]  (.SI(n74), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.QN(n50), 
	.Q(n167), 
	.D(n130), 
	.CK(CLK));
   OAI22X2M U33 (.Y(FUN[2]), 
	.B1(n119), 
	.B0(n45), 
	.A1(n118), 
	.A0(n48));
   NOR2X3M U35 (.Y(Addr[2]), 
	.B(n45), 
	.A(n121));
   NAND4X2M U36 (.Y(n98), 
	.D(n72), 
	.C(n101), 
	.B(n150), 
	.A(enable_pulse));
   OAI22X1M U37 (.Y(FUN[0]), 
	.B1(n119), 
	.B0(n47), 
	.A1(n118), 
	.A0(n51));
   OAI22X1M U38 (.Y(FUN[1]), 
	.B1(n119), 
	.B0(n46), 
	.A1(n118), 
	.A0(n49));
   INVX2M U39 (.Y(n34), 
	.A(n76));
   NAND3BX2M U40 (.Y(n76), 
	.C(n71), 
	.B(n82), 
	.AN(FIFO_FULL));
   INVX2M U41 (.Y(n53), 
	.A(n78));
   INVX2M U42 (.Y(n52), 
	.A(n100));
   INVX2M U43 (.Y(n70), 
	.A(n79));
   NAND2BX2M U44 (.Y(n118), 
	.B(ALU_En), 
	.AN(n116));
   NAND2X2M U45 (.Y(n119), 
	.B(ALU_En), 
	.A(n66));
   NOR2BX2M U46 (.Y(n121), 
	.B(Rd_En), 
	.AN(n102));
   NOR3X2M U47 (.Y(n108), 
	.C(n89), 
	.B(FIFO_FULL), 
	.A(n105));
   NAND3X2M U48 (.Y(n79), 
	.C(n104), 
	.B(n72), 
	.A(n150));
   OAI21BX1M U49 (.Y(WR_INC), 
	.B0N(n106), 
	.A1(n105), 
	.A0(FIFO_FULL));
   NOR4X1M U50 (.Y(n106), 
	.D(n73), 
	.C(n150), 
	.B(n72), 
	.A(n68));
   NAND2X2M U51 (.Y(n80), 
	.B(n104), 
	.A(n103));
   NAND4X2M U52 (.Y(n116), 
	.D(n147), 
	.C(n57), 
	.B(n120), 
	.A(n88));
   NAND2X2M U53 (.Y(n82), 
	.B(n117), 
	.A(n116));
   NAND3X2M U54 (.Y(Wr_En), 
	.C(n102), 
	.B(n79), 
	.A(n80));
   INVX2M U55 (.Y(n71), 
	.A(n105));
   AOI221XLM U56 (.Y(n83), 
	.C0(Rd_En), 
	.B1(n67), 
	.B0(n78), 
	.A1(n71), 
	.A0(n89));
   INVX2M U57 (.Y(n67), 
	.A(n89));
   OAI22X1M U58 (.Y(n136), 
	.B1(n149), 
	.B0(n56), 
	.A1(n98), 
	.A0(n49));
   OAI22X1M U59 (.Y(n135), 
	.B1(n148), 
	.B0(n56), 
	.A1(n98), 
	.A0(n48));
   OAI22X1M U60 (.Y(n133), 
	.B1(n147), 
	.B0(n56), 
	.A1(n98), 
	.A0(n38));
   OAI22X1M U61 (.Y(n132), 
	.B1(n146), 
	.B0(n56), 
	.A1(n98), 
	.A0(n37));
   OAI22X1M U62 (.Y(n131), 
	.B1(n74), 
	.B0(n56), 
	.A1(n98), 
	.A0(n36));
   OAI22X1M U63 (.Y(n145), 
	.B1(n57), 
	.B0(n56), 
	.A1(n98), 
	.A0(n51));
   INVX2M U64 (.Y(n56), 
	.A(n98));
   NAND3X2M U65 (.Y(n99), 
	.C(n103), 
	.B(n68), 
	.A(n73));
   NOR2X2M U67 (.Y(n78), 
	.B(n55), 
	.A(n99));
   NOR2X2M U69 (.Y(n100), 
	.B(n55), 
	.A(n80));
   INVX2M U70 (.Y(ALU_En), 
	.A(n75));
   NAND4X2M U71 (.Y(next_state[2]), 
	.D(n81), 
	.C(n80), 
	.B(n79), 
	.A(n75));
   AOI21BX2M U72 (.Y(n81), 
	.B0N(n83), 
	.A1(n82), 
	.A0(n78));
   INVX2M U73 (.Y(n66), 
	.A(n117));
   OAI211X2M U74 (.Y(Gate_En), 
	.C0(n79), 
	.B0(n75), 
	.A1(n117), 
	.A0(n99));
   NOR2X2M U75 (.Y(n104), 
	.B(current_state[3]), 
	.A(n73));
   AND3X2M U76 (.Y(Rd_En), 
	.C(current_state[1]), 
	.B(n150), 
	.A(n104));
   INVX2M U77 (.Y(n73), 
	.A(current_state[2]));
   OAI21X2M U78 (.Y(Addr[0]), 
	.B0(n79), 
	.A1(n47), 
	.A0(n121));
   NOR2X4M U79 (.Y(Addr[3]), 
	.B(n44), 
	.A(n121));
   NOR4X1M U80 (.Y(n120), 
	.D(Stored_Frame1[5]), 
	.C(Stored_Frame1[1]), 
	.B(n148), 
	.A(n74));
   OAI222X1M U81 (.Y(Wr_D[1]), 
	.C1(n102), 
	.C0(n49), 
	.B1(n64), 
	.B0(n79), 
	.A1(n46), 
	.A0(n80));
   OAI222X1M U82 (.Y(Wr_D[2]), 
	.C1(n102), 
	.C0(n48), 
	.B1(n63), 
	.B0(n79), 
	.A1(n45), 
	.A0(n80));
   OAI222X1M U83 (.Y(Wr_D[3]), 
	.C1(n102), 
	.C0(n39), 
	.B1(n62), 
	.B0(n79), 
	.A1(n44), 
	.A0(n80));
   OAI222X1M U84 (.Y(Wr_D[0]), 
	.C1(n102), 
	.C0(n51), 
	.B1(n65), 
	.B0(n79), 
	.A1(n47), 
	.A0(n80));
   OAI222X1M U85 (.Y(Wr_D[4]), 
	.C1(n102), 
	.C0(n38), 
	.B1(n61), 
	.B0(n79), 
	.A1(n43), 
	.A0(n80));
   OAI222X1M U86 (.Y(Wr_D[5]), 
	.C1(n102), 
	.C0(n37), 
	.B1(n60), 
	.B0(n79), 
	.A1(n42), 
	.A0(n80));
   OAI222X1M U87 (.Y(Wr_D[6]), 
	.C1(n102), 
	.C0(n36), 
	.B1(n59), 
	.B0(n79), 
	.A1(n41), 
	.A0(n80));
   OAI222X1M U88 (.Y(Wr_D[7]), 
	.C1(n102), 
	.C0(n35), 
	.B1(n58), 
	.B0(n79), 
	.A1(n40), 
	.A0(n80));
   NOR4X1M U89 (.Y(n85), 
	.D(Stored_Frame1[6]), 
	.C(Stored_Frame1[2]), 
	.B(n149), 
	.A(n146));
   NOR2X2M U90 (.Y(n103), 
	.B(current_state[1]), 
	.A(n150));
   NAND4X2M U91 (.Y(n102), 
	.D(n68), 
	.C(n73), 
	.B(n150), 
	.A(current_state[1]));
   NAND4X2M U92 (.Y(n89), 
	.D(Stored_Frame1[0]), 
	.C(Stored_Frame1[4]), 
	.B(n88), 
	.A(n85));
   NAND4X2M U93 (.Y(n117), 
	.D(n120), 
	.C(Stored_Frame1[0]), 
	.B(Stored_Frame1[4]), 
	.A(n88));
   INVX2M U94 (.Y(n150), 
	.A(current_state[0]));
   NAND3X2M U95 (.Y(n105), 
	.C(current_state[1]), 
	.B(n104), 
	.A(current_state[0]));
   INVX2M U96 (.Y(n72), 
	.A(current_state[1]));
   OAI2BB1X2M U97 (.Y(WR_DATA[0]), 
	.B0(n115), 
	.A1N(n106), 
	.A0N(ALU_OUT[8]));
   AOI22X1M U98 (.Y(n115), 
	.B1(n108), 
	.B0(Rd_D[0]), 
	.A1(n34), 
	.A0(ALU_OUT[0]));
   OAI2BB1X2M U99 (.Y(WR_DATA[1]), 
	.B0(n114), 
	.A1N(n106), 
	.A0N(ALU_OUT[9]));
   AOI22X1M U100 (.Y(n114), 
	.B1(n108), 
	.B0(Rd_D[1]), 
	.A1(n34), 
	.A0(ALU_OUT[1]));
   OAI2BB1X2M U101 (.Y(WR_DATA[2]), 
	.B0(n113), 
	.A1N(n106), 
	.A0N(ALU_OUT[10]));
   AOI22X1M U102 (.Y(n113), 
	.B1(n108), 
	.B0(Rd_D[2]), 
	.A1(n34), 
	.A0(ALU_OUT[2]));
   OAI2BB1X2M U103 (.Y(WR_DATA[3]), 
	.B0(n112), 
	.A1N(n106), 
	.A0N(ALU_OUT[11]));
   AOI22X1M U104 (.Y(n112), 
	.B1(n108), 
	.B0(Rd_D[3]), 
	.A1(n34), 
	.A0(ALU_OUT[3]));
   OAI2BB1X2M U105 (.Y(WR_DATA[4]), 
	.B0(n111), 
	.A1N(n106), 
	.A0N(ALU_OUT[12]));
   AOI22X1M U106 (.Y(n111), 
	.B1(n108), 
	.B0(Rd_D[4]), 
	.A1(n34), 
	.A0(ALU_OUT[4]));
   OAI2BB1X2M U107 (.Y(WR_DATA[5]), 
	.B0(n110), 
	.A1N(n106), 
	.A0N(ALU_OUT[13]));
   AOI22X1M U108 (.Y(n110), 
	.B1(n108), 
	.B0(Rd_D[5]), 
	.A1(n34), 
	.A0(ALU_OUT[5]));
   OAI2BB1X2M U109 (.Y(WR_DATA[6]), 
	.B0(n109), 
	.A1N(n106), 
	.A0N(ALU_OUT[14]));
   AOI22X1M U110 (.Y(n109), 
	.B1(n108), 
	.B0(Rd_D[6]), 
	.A1(n34), 
	.A0(ALU_OUT[6]));
   OAI2BB1X2M U111 (.Y(WR_DATA[7]), 
	.B0(n107), 
	.A1N(n106), 
	.A0N(ALU_OUT[15]));
   AOI22X1M U112 (.Y(n107), 
	.B1(n108), 
	.B0(Rd_D[7]), 
	.A1(n34), 
	.A0(ALU_OUT[7]));
   INVX2M U113 (.Y(n68), 
	.A(current_state[3]));
   NOR2X2M U114 (.Y(Addr[1]), 
	.B(n46), 
	.A(n121));
   INVX2M U115 (.Y(n148), 
	.A(Stored_Frame1[2]));
   INVX2M U116 (.Y(n149), 
	.A(Stored_Frame1[1]));
   INVX2M U117 (.Y(n74), 
	.A(Stored_Frame1[6]));
   INVX2M U118 (.Y(n146), 
	.A(Stored_Frame1[5]));
   AOI222X1M U119 (.Y(n93), 
	.C1(n70), 
	.C0(enable_pulse), 
	.B1(n89), 
	.B0(n71), 
	.A1(Rd_En), 
	.A0(Rd_D_Valid));
   AOI211X2M U120 (.Y(n95), 
	.C0(n98), 
	.B0(n39), 
	.A1(n97), 
	.A0(n96));
   NAND4X2M U121 (.Y(n96), 
	.D(n36), 
	.C(n48), 
	.B(Sync_Frame[1]), 
	.A(Sync_Frame[5]));
   NAND4X2M U122 (.Y(n97), 
	.D(n37), 
	.C(n49), 
	.B(Sync_Frame[2]), 
	.A(Sync_Frame[6]));
   NOR2X2M U123 (.Y(n88), 
	.B(n54), 
	.A(n50));
   NOR4X1M U124 (.Y(n87), 
	.D(current_state[3]), 
	.C(current_state[2]), 
	.B(n150), 
	.A(n72));
   NAND3X2M U125 (.Y(n75), 
	.C(current_state[3]), 
	.B(current_state[2]), 
	.A(n103));
   XNOR2X2M U126 (.Y(n94), 
	.B(Sync_Frame[0]), 
	.A(Sync_Frame[4]));
   OAI22X1M U127 (.Y(n134), 
	.B1(n54), 
	.B0(n56), 
	.A1(n39), 
	.A0(n98));
   OAI22X1M U128 (.Y(n130), 
	.B1(n50), 
	.B0(n56), 
	.A1(n35), 
	.A0(n98));
   OAI22X1M U129 (.Y(n122), 
	.B1(n65), 
	.B0(n100), 
	.A1(n52), 
	.A0(n51));
   OAI22X1M U130 (.Y(n123), 
	.B1(n64), 
	.B0(n100), 
	.A1(n52), 
	.A0(n49));
   OAI22X1M U131 (.Y(n124), 
	.B1(n63), 
	.B0(n100), 
	.A1(n52), 
	.A0(n48));
   OAI22X1M U132 (.Y(n125), 
	.B1(n62), 
	.B0(n100), 
	.A1(n52), 
	.A0(n39));
   OAI22X1M U133 (.Y(n126), 
	.B1(n61), 
	.B0(n100), 
	.A1(n52), 
	.A0(n38));
   OAI22X1M U134 (.Y(n127), 
	.B1(n60), 
	.B0(n100), 
	.A1(n52), 
	.A0(n37));
   OAI22X1M U135 (.Y(n128), 
	.B1(n59), 
	.B0(n100), 
	.A1(n52), 
	.A0(n36));
   OAI22X1M U136 (.Y(n129), 
	.B1(n58), 
	.B0(n100), 
	.A1(n52), 
	.A0(n35));
   OAI22X1M U137 (.Y(n140), 
	.B1(n43), 
	.B0(n78), 
	.A1(n38), 
	.A0(n53));
   OAI22X1M U138 (.Y(n139), 
	.B1(n42), 
	.B0(n78), 
	.A1(n37), 
	.A0(n53));
   OAI22X1M U139 (.Y(n138), 
	.B1(n41), 
	.B0(n78), 
	.A1(n36), 
	.A0(n53));
   OAI22X1M U140 (.Y(n137), 
	.B1(n40), 
	.B0(n78), 
	.A1(n35), 
	.A0(n53));
   OAI22X1M U141 (.Y(n144), 
	.B1(n47), 
	.B0(n78), 
	.A1(n51), 
	.A0(n53));
   OAI22X1M U142 (.Y(n143), 
	.B1(n46), 
	.B0(n78), 
	.A1(n49), 
	.A0(n53));
   OAI22X1M U143 (.Y(n142), 
	.B1(n45), 
	.B0(n78), 
	.A1(n48), 
	.A0(n53));
   OAI22X1M U144 (.Y(n141), 
	.B1(n44), 
	.B0(n78), 
	.A1(n39), 
	.A0(n53));
   OAI2B11X2M U145 (.Y(next_state[1]), 
	.C0(n84), 
	.B0(n83), 
	.A1N(OUT_Valid), 
	.A0(n75));
   AOI31X2M U146 (.Y(n84), 
	.B0(n87), 
	.A2(n86), 
	.A1(n78), 
	.A0(n85));
   AND3X2M U147 (.Y(n86), 
	.C(n57), 
	.B(n147), 
	.A(n88));
   OAI211X2M U148 (.Y(next_state[3]), 
	.C0(n77), 
	.B0(n76), 
	.A1(n75), 
	.A0(OUT_Valid));
   AOI22X1M U149 (.Y(n77), 
	.B1(n66), 
	.B0(n78), 
	.A1(n70), 
	.A0(enable_pulse));
   NOR2X2M U150 (.Y(n101), 
	.B(current_state[2]), 
	.A(current_state[3]));
   NAND4X2M U151 (.Y(next_state[0]), 
	.D(n93), 
	.C(n92), 
	.B(n91), 
	.A(n90));
   OAI21BX1M U152 (.Y(n90), 
	.B0N(n99), 
	.A1(n89), 
	.A0(n55));
   OAI2B1X2M U153 (.Y(n91), 
	.B0(n55), 
	.A1N(n80), 
	.A0(n87));
   AOI31X2M U154 (.Y(n92), 
	.B0(ALU_En), 
	.A2(n95), 
	.A1(Sync_Frame[7]), 
	.A0(n94));
   INVX2M U155 (.Y(n49), 
	.A(Sync_Frame[1]));
   INVX2M U156 (.Y(n48), 
	.A(Sync_Frame[2]));
   INVX2M U157 (.Y(n55), 
	.A(enable_pulse));
   INVX2M U158 (.Y(n37), 
	.A(Sync_Frame[5]));
   INVX2M U159 (.Y(n36), 
	.A(Sync_Frame[6]));
   INVX2M U160 (.Y(n39), 
	.A(Sync_Frame[3]));
   INVX2M U161 (.Y(n51), 
	.A(Sync_Frame[0]));
   INVX2M U162 (.Y(n57), 
	.A(Stored_Frame1[0]));
   INVX2M U163 (.Y(n147), 
	.A(Stored_Frame1[4]));
   INVX2M U164 (.Y(n38), 
	.A(Sync_Frame[4]));
   INVX2M U165 (.Y(n35), 
	.A(Sync_Frame[7]));
   OAI22X2M U166 (.Y(FUN[3]), 
	.B1(n119), 
	.B0(n44), 
	.A1(n118), 
	.A0(n39));
   INVX2M U3 (.Y(CLK_DIV_EN), 
	.A(LTIE_LTIELO_NET));
endmodule

module Integer_ClkDiv_ratio_Width8_DW01_inc_0 (
	A, 
	SUM);
   input [6:0] A;
   output [6:0] SUM;

   // Internal wires
   wire [6:2] carry;

   ADDHX1M U1_1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.B(carry[5]), 
	.A(A[5]));
   ADDHX1M U1_1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.B(carry[4]), 
	.A(A[4]));
   ADDHX1M U1_1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.B(A[0]), 
	.A(A[1]));
   ADDHX1M U1_1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.B(carry[3]), 
	.A(A[3]));
   ADDHX1M U1_1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.B(carry[2]), 
	.A(A[2]));
   CLKXOR2X2M U1 (.Y(SUM[6]), 
	.B(A[6]), 
	.A(carry[6]));
   CLKINVX1M U2 (.Y(SUM[0]), 
	.A(A[0]));
endmodule

module Integer_ClkDiv_ratio_Width8_test_1 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	UART_CLK_M__L1_N0, 
	UART_CLK_M__L6_N1);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input UART_CLK_M__L1_N0;
   input UART_CLK_M__L6_N1;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire N0;
   wire New_clk;
   wire Flag;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire N44;
   wire N45;
   wire n17;
   wire n29;
   wire n30;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n16;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire [6:0] Half_Div;
   wire [6:0] Count;

//   assign test_so = New_clk ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   SDFFSX1M New_clk_reg (.SN(i_rst_n), 
	.SI(Flag), 
	.SE(test_se), 
	.QN(n17), 
	.Q(test_so), 
	.D(n30), 
	.CK(UART_CLK_M__L1_N0));
   SDFFRQX2M Flag_reg (.SI(n41), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Flag), 
	.D(n29), 
	.CK(i_ref_clk));
   SDFFRQX2M \Count_reg[6]  (.SI(Count[5]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Count[6]), 
	.D(N45), 
	.CK(i_ref_clk));
   SDFFRQX2M \Count_reg[5]  (.SI(Count[4]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Count[5]), 
	.D(N44), 
	.CK(i_ref_clk));
   SDFFRQX2M \Count_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Count[0]), 
	.D(N39), 
	.CK(i_ref_clk));
   SDFFRQX2M \Count_reg[4]  (.SI(n56), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Count[4]), 
	.D(N43), 
	.CK(i_ref_clk));
   SDFFRQX2M \Count_reg[1]  (.SI(Count[0]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Count[1]), 
	.D(N40), 
	.CK(i_ref_clk));
   SDFFRQX2M \Count_reg[3]  (.SI(Count[2]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Count[3]), 
	.D(N42), 
	.CK(i_ref_clk));
   SDFFRQX2M \Count_reg[2]  (.SI(Count[1]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Count[2]), 
	.D(N41), 
	.CK(i_ref_clk));
   AOI21BX2M U5 (.Y(n1), 
	.B0N(n3), 
	.A1(i_div_ratio[3]), 
	.A0(n2));
   OR2X2M U6 (.Y(n2), 
	.B(i_div_ratio[1]), 
	.A(i_div_ratio[2]));
   INVX2M U14 (.Y(n16), 
	.A(i_div_ratio[5]));
   MX2X2M U15 (.Y(o_div_clk), 
	.S0(N0), 
	.B(test_so), 
	.A(UART_CLK_M__L6_N1));
   CLKINVX1M U16 (.Y(Half_Div[0]), 
	.A(i_div_ratio[1]));
   OAI2BB1X1M U17 (.Y(Half_Div[1]), 
	.B0(n2), 
	.A1N(i_div_ratio[2]), 
	.A0N(i_div_ratio[1]));
   OR2X1M U18 (.Y(n3), 
	.B(i_div_ratio[3]), 
	.A(n2));
   NOR2X1M U19 (.Y(n4), 
	.B(i_div_ratio[4]), 
	.A(n3));
   AO21XLM U20 (.Y(Half_Div[3]), 
	.B0(n4), 
	.A1(i_div_ratio[4]), 
	.A0(n3));
   CLKNAND2X2M U21 (.Y(n5), 
	.B(n16), 
	.A(n4));
   OAI21X1M U22 (.Y(Half_Div[4]), 
	.B0(n5), 
	.A1(n16), 
	.A0(n4));
   XNOR2X1M U23 (.Y(Half_Div[5]), 
	.B(n5), 
	.A(i_div_ratio[6]));
   NOR2X1M U24 (.Y(n6), 
	.B(n5), 
	.A(i_div_ratio[6]));
   CLKXOR2X2M U25 (.Y(Half_Div[6]), 
	.B(n6), 
	.A(i_div_ratio[7]));
   MXI2X1M U26 (.Y(n30), 
	.S0(n19), 
	.B(n18), 
	.A(n17));
   NOR2X1M U27 (.Y(n18), 
	.B(n20), 
	.A(n17));
   NOR2X1M U28 (.Y(n29), 
	.B(n21), 
	.A(n20));
   MXI2X1M U29 (.Y(n21), 
	.S0(Flag), 
	.B(n23), 
	.A(n22));
   NOR2X1M U30 (.Y(n23), 
	.B(n24), 
	.A(n22));
   CLKINVX1M U31 (.Y(n22), 
	.A(n25));
   NOR2BX1M U32 (.Y(N45), 
	.B(n19), 
	.AN(N24));
   NOR2BX1M U33 (.Y(N44), 
	.B(n19), 
	.AN(N23));
   NOR2BX1M U34 (.Y(N43), 
	.B(n19), 
	.AN(N22));
   NOR2BX1M U35 (.Y(N42), 
	.B(n19), 
	.AN(N21));
   NOR2BX1M U36 (.Y(N41), 
	.B(n19), 
	.AN(N20));
   NOR2BX1M U37 (.Y(N40), 
	.B(n19), 
	.AN(N19));
   NOR2BX1M U38 (.Y(N39), 
	.B(n19), 
	.AN(N18));
   OAI211X1M U39 (.Y(n19), 
	.C0(n27), 
	.B0(n25), 
	.A1(n26), 
	.A0(i_div_ratio[0]));
   NOR2X1M U40 (.Y(n27), 
	.B(n20), 
	.A(n24));
   CLKNAND2X2M U41 (.Y(n25), 
	.B(i_div_ratio[0]), 
	.A(n28));
   MXI2X1M U42 (.Y(n28), 
	.S0(Flag), 
	.B(n31), 
	.A(n26));
   NAND4X1M U43 (.Y(n31), 
	.D(n35), 
	.C(n34), 
	.B(n33), 
	.A(n32));
   NOR4X1M U44 (.Y(n35), 
	.D(n39), 
	.C(n38), 
	.B(n37), 
	.A(n36));
   CLKXOR2X2M U45 (.Y(n39), 
	.B(Count[3]), 
	.A(i_div_ratio[4]));
   CLKXOR2X2M U46 (.Y(n38), 
	.B(Count[2]), 
	.A(i_div_ratio[3]));
   CLKXOR2X2M U47 (.Y(n37), 
	.B(Count[1]), 
	.A(i_div_ratio[2]));
   CLKXOR2X2M U48 (.Y(n36), 
	.B(Count[0]), 
	.A(i_div_ratio[1]));
   CLKXOR2X2M U49 (.Y(n34), 
	.B(i_div_ratio[6]), 
	.A(n40));
   CLKXOR2X2M U50 (.Y(n33), 
	.B(i_div_ratio[7]), 
	.A(n41));
   CLKXOR2X2M U51 (.Y(n32), 
	.B(i_div_ratio[5]), 
	.A(n42));
   NAND4BX1M U52 (.Y(n26), 
	.D(n45), 
	.C(n44), 
	.B(n43), 
	.AN(n24));
   NOR4X1M U53 (.Y(n45), 
	.D(n49), 
	.C(n48), 
	.B(n47), 
	.A(n46));
   AOI21X1M U54 (.Y(n44), 
	.B0(n51), 
	.A1(n50), 
	.A0(Half_Div[0]));
   CLKNAND2X2M U55 (.Y(n43), 
	.B(n52), 
	.A(Half_Div[1]));
   OAI32X1M U56 (.Y(n24), 
	.B1(n41), 
	.B0(Half_Div[6]), 
	.A2(n49), 
	.A1(n48), 
	.A0(n53));
   CLKINVX1M U57 (.Y(n41), 
	.A(Count[6]));
   NOR2BX1M U58 (.Y(n49), 
	.B(Count[5]), 
	.AN(Half_Div[5]));
   NOR2BX1M U59 (.Y(n48), 
	.B(Count[6]), 
	.AN(Half_Div[6]));
   CLKINVX1M U60 (.Y(n53), 
	.A(n54));
   OAI222X1M U61 (.Y(n54), 
	.C1(Half_Div[4]), 
	.C0(n42), 
	.B1(n46), 
	.B0(n55), 
	.A1(Half_Div[5]), 
	.A0(n40));
   AND2X1M U62 (.Y(n46), 
	.B(n42), 
	.A(Half_Div[4]));
   CLKINVX1M U63 (.Y(n42), 
	.A(Count[4]));
   OA22X1M U64 (.Y(n55), 
	.B1(n57), 
	.B0(n51), 
	.A1(n56), 
	.A0(Half_Div[3]));
   AOI32X1M U65 (.Y(n57), 
	.B1(n1), 
	.B0(Count[2]), 
	.A2(n60), 
	.A1(n59), 
	.A0(n58));
   OAI21X1M U66 (.Y(n60), 
	.B0(n52), 
	.A1(n50), 
	.A0(Half_Div[0]));
   CLKINVX1M U67 (.Y(n59), 
	.A(n47));
   NOR2X1M U68 (.Y(n47), 
	.B(Count[2]), 
	.A(n1));
   OAI31X1M U69 (.Y(n58), 
	.B0(Half_Div[1]), 
	.A2(n50), 
	.A1(Half_Div[0]), 
	.A0(n52));
   CLKINVX1M U70 (.Y(n50), 
	.A(Count[0]));
   CLKINVX1M U71 (.Y(n52), 
	.A(Count[1]));
   NOR2BX1M U72 (.Y(n51), 
	.B(Count[3]), 
	.AN(Half_Div[3]));
   CLKINVX1M U73 (.Y(n56), 
	.A(Count[3]));
   CLKINVX1M U74 (.Y(n40), 
	.A(Count[5]));
   CLKINVX1M U75 (.Y(N0), 
	.A(n20));
   OAI21X1M U76 (.Y(n20), 
	.B0(HTIE_LTIEHI_NET), 
	.A1(n62), 
	.A0(n61));
   OR3X1M U77 (.Y(n62), 
	.C(i_div_ratio[1]), 
	.B(i_div_ratio[3]), 
	.A(i_div_ratio[2]));
   OR4X1M U78 (.Y(n61), 
	.D(i_div_ratio[7]), 
	.C(i_div_ratio[6]), 
	.B(i_div_ratio[5]), 
	.A(i_div_ratio[4]));
   Integer_ClkDiv_ratio_Width8_DW01_inc_0 add_73 (.A({ Count[6],
		Count[5],
		Count[4],
		Count[3],
		Count[2],
		Count[1],
		Count[0] }), 
	.SUM({ N24,
		N23,
		N22,
		N21,
		N20,
		N19,
		N18 }));
endmodule

module Integer_ClkDiv_ratio_Width4_test_1 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	UART_CLK_M__L2_N1, 
	UART_CLK_M__L7_N0);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [3:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input UART_CLK_M__L2_N1;
   input UART_CLK_M__L7_N0;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire N0;
   wire New_clk;
   wire N31;
   wire N32;
   wire N33;
   wire n12;
   wire n13;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire [2:0] Count;

//   assign test_so = New_clk ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   SDFFRX1M Flag_reg (.SI(n5), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.QN(n12), 
	.Q(n6), 
	.D(n33), 
	.CK(i_ref_clk));
   SDFFRQX2M \Count_reg[2]  (.SI(n4), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Count[2]), 
	.D(N33), 
	.CK(i_ref_clk));
   SDFFRQX2M \Count_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Count[0]), 
	.D(N31), 
	.CK(i_ref_clk));
   SDFFRQX2M \Count_reg[1]  (.SI(n3), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Count[1]), 
	.D(N32), 
	.CK(i_ref_clk));
   SDFFSX1M New_clk_reg (.SN(i_rst_n), 
	.SI(n6), 
	.SE(test_se), 
	.QN(n13), 
	.Q(test_so), 
	.D(n34), 
	.CK(UART_CLK_M__L2_N1));
   OAI32X1M U9 (.Y(n18), 
	.B1(n5), 
	.B0(n31), 
	.A2(n30), 
	.A1(n28), 
	.A0(n29));
   OAI2B11X2M U10 (.Y(n21), 
	.C0(n25), 
	.B0(n20), 
	.A1N(n24), 
	.A0(i_div_ratio[0]));
   NOR2X2M U11 (.Y(n25), 
	.B(n19), 
	.A(n18));
   AOI21BX2M U12 (.Y(n27), 
	.B0N(n32), 
	.A1(i_div_ratio[2]), 
	.A0(i_div_ratio[1]));
   OR2X2M U13 (.Y(n32), 
	.B(i_div_ratio[1]), 
	.A(i_div_ratio[2]));
   AND2X2M U14 (.Y(n31), 
	.B(n32), 
	.A(i_div_ratio[3]));
   INVX2M U15 (.Y(N0), 
	.A(n19));
   NOR2X2M U16 (.Y(n29), 
	.B(n27), 
	.A(Count[1]));
   AOI22X1M U17 (.Y(n30), 
	.B1(i_div_ratio[1]), 
	.B0(Count[0]), 
	.A1(n27), 
	.A0(Count[1]));
   AOI211X2M U18 (.Y(n24), 
	.C0(n26), 
	.B0(n18), 
	.A1(n3), 
	.A0(n2));
   INVX2M U19 (.Y(n2), 
	.A(i_div_ratio[1]));
   OAI21BX1M U20 (.Y(n26), 
	.B0N(n28), 
	.A1(Count[1]), 
	.A0(n27));
   OAI32X1M U21 (.Y(N33), 
	.B1(n21), 
	.B0(n5), 
	.A2(n3), 
	.A1(n4), 
	.A0(n21));
   INVX2M U22 (.Y(n4), 
	.A(Count[1]));
   OAI21X2M U23 (.Y(n34), 
	.B0(n22), 
	.A1(n21), 
	.A0(n13));
   OAI21X2M U24 (.Y(n22), 
	.B0(n21), 
	.A1(n13), 
	.A0(n19));
   NAND3X2M U25 (.Y(n20), 
	.C(i_div_ratio[0]), 
	.B(n12), 
	.A(n24));
   NOR2X2M U26 (.Y(N32), 
	.B(n21), 
	.A(n23));
   CLKXOR2X2M U27 (.Y(n23), 
	.B(Count[1]), 
	.A(n3));
   NOR2X2M U28 (.Y(N31), 
	.B(n21), 
	.A(Count[0]));
   NOR2BX2M U29 (.Y(n28), 
	.B(Count[2]), 
	.AN(n31));
   OAI21X2M U30 (.Y(n19), 
	.B0(HTIE_LTIEHI_NET), 
	.A1(n32), 
	.A0(i_div_ratio[3]));
   OAI32X1M U31 (.Y(n33), 
	.B1(n19), 
	.B0(n20), 
	.A2(n19), 
	.A1(n18), 
	.A0(n12));
   INVX2M U32 (.Y(n3), 
	.A(Count[0]));
   INVX2M U33 (.Y(n5), 
	.A(Count[2]));
   MX2X2M U34 (.Y(o_div_clk), 
	.S0(N0), 
	.B(test_so), 
	.A(UART_CLK_M__L7_N0));
endmodule

module RX_CLKDIV_MUX_Width4 (
	Input, 
	MUX_Out);
   input [5:0] Input;
   output [3:0] MUX_Out;

   // Internal wires
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n1;
   wire n2;
   wire n3;
   wire n4;

   NAND4BX1M U3 (.Y(n6), 
	.D(n1), 
	.C(n2), 
	.B(Input[3]), 
	.AN(Input[4]));
   NAND4BX1M U4 (.Y(n7), 
	.D(n1), 
	.C(n2), 
	.B(Input[4]), 
	.AN(Input[3]));
   NOR3X2M U5 (.Y(MUX_Out[1]), 
	.C(Input[0]), 
	.B(Input[1]), 
	.A(n7));
   NOR4X1M U6 (.Y(MUX_Out[3]), 
	.D(Input[4]), 
	.C(Input[5]), 
	.B(Input[3]), 
	.A(n5));
   NAND3X2M U7 (.Y(n5), 
	.C(Input[2]), 
	.B(n3), 
	.A(n4));
   NOR3X2M U8 (.Y(MUX_Out[2]), 
	.C(Input[0]), 
	.B(Input[1]), 
	.A(n6));
   INVX2M U9 (.Y(n2), 
	.A(Input[2]));
   INVX2M U10 (.Y(n4), 
	.A(Input[0]));
   INVX2M U11 (.Y(n3), 
	.A(Input[1]));
   INVX2M U12 (.Y(n1), 
	.A(Input[5]));
   OAI211X2M U13 (.Y(MUX_Out[0]), 
	.C0(n3), 
	.B0(n4), 
	.A1(n9), 
	.A0(n8));
   NOR4X1M U14 (.Y(n8), 
	.D(n2), 
	.C(Input[3]), 
	.B(Input[4]), 
	.A(Input[5]));
   NAND2X2M U15 (.Y(n9), 
	.B(n6), 
	.A(n7));
endmodule

module Data_Sampling_test_1 (
	CLK, 
	RST, 
	En, 
	Prescale, 
	RX_In, 
	Edge_Count, 
	Sampeld_Bit, 
	test_si, 
	test_so, 
	test_se, 
	RX_CLK_M__L3_N1);
   input CLK;
   input RST;
   input En;
   input [5:0] Prescale;
   input RX_In;
   input [5:0] Edge_Count;
   output Sampeld_Bit;
   input test_si;
   output test_so;
   input test_se;
   input RX_CLK_M__L3_N1;

   // Internal wires
   wire N25;
   wire n23;
   wire n24;
   wire n25;
   wire \add_28/carry[4] ;
   wire \add_28/carry[3] ;
   wire \add_28/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire [4:0] Middle_Sample_Plus;
   wire [4:0] Middle_Sample_minus;
   wire [2:0] Samples;

   assign test_so = Samples[2] ;

   SDFFRQX2M \Samples_reg[2]  (.SI(Samples[1]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Samples[2]), 
	.D(n25), 
	.CK(CLK));
   SDFFRQX2M \Samples_reg[1]  (.SI(Samples[0]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Samples[1]), 
	.D(n24), 
	.CK(RX_CLK_M__L3_N1));
   SDFFRQX2M \Samples_reg[0]  (.SI(Sampeld_Bit), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Samples[0]), 
	.D(n23), 
	.CK(RX_CLK_M__L3_N1));
   SDFFRQX2M Sampeld_Bit_reg (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Sampeld_Bit), 
	.D(N25), 
	.CK(CLK));
   INVX2M U4 (.Y(n4), 
	.A(Prescale[3]));
   ADDHX1M U5 (.S(Middle_Sample_Plus[2]), 
	.CO(\add_28/carry[3] ), 
	.B(\add_28/carry[2] ), 
	.A(Prescale[3]));
   ADDHX1M U6 (.S(Middle_Sample_Plus[1]), 
	.CO(\add_28/carry[2] ), 
	.B(Prescale[1]), 
	.A(Prescale[2]));
   ADDHX1M U10 (.S(Middle_Sample_Plus[3]), 
	.CO(\add_28/carry[4] ), 
	.B(\add_28/carry[3] ), 
	.A(Prescale[4]));
   CLKXOR2X2M U11 (.Y(Middle_Sample_Plus[4]), 
	.B(Prescale[5]), 
	.A(\add_28/carry[4] ));
   CLKINVX1M U12 (.Y(Middle_Sample_minus[0]), 
	.A(Prescale[1]));
   NOR2X1M U13 (.Y(n1), 
	.B(Prescale[1]), 
	.A(Prescale[2]));
   AO21XLM U14 (.Y(Middle_Sample_minus[1]), 
	.B0(n1), 
	.A1(Prescale[2]), 
	.A0(Prescale[1]));
   CLKNAND2X2M U15 (.Y(n2), 
	.B(n4), 
	.A(n1));
   OAI21X1M U16 (.Y(Middle_Sample_minus[2]), 
	.B0(n2), 
	.A1(n4), 
	.A0(n1));
   XNOR2X1M U17 (.Y(Middle_Sample_minus[3]), 
	.B(n2), 
	.A(Prescale[4]));
   NOR2X1M U18 (.Y(n3), 
	.B(n2), 
	.A(Prescale[4]));
   CLKXOR2X2M U19 (.Y(Middle_Sample_minus[4]), 
	.B(n3), 
	.A(Prescale[5]));
   MXI2X1M U20 (.Y(n25), 
	.S0(n11), 
	.B(n6), 
	.A(n5));
   NOR2X1M U21 (.Y(n11), 
	.B(n13), 
	.A(n12));
   NAND4X1M U22 (.Y(n13), 
	.D(n17), 
	.C(n16), 
	.B(n15), 
	.A(n14));
   CLKXOR2X2M U23 (.Y(n17), 
	.B(Middle_Sample_Plus[1]), 
	.A(n18));
   XNOR2X1M U24 (.Y(n16), 
	.B(Middle_Sample_Plus[2]), 
	.A(Edge_Count[2]));
   XNOR2X1M U25 (.Y(n15), 
	.B(Middle_Sample_Plus[3]), 
	.A(Edge_Count[3]));
   CLKXOR2X2M U26 (.Y(n14), 
	.B(Middle_Sample_Plus[4]), 
	.A(n19));
   NAND4BX1M U27 (.Y(n12), 
	.D(n22), 
	.C(n21), 
	.B(n20), 
	.AN(Edge_Count[5]));
   XNOR2X1M U28 (.Y(n20), 
	.B(Middle_Sample_minus[0]), 
	.A(Edge_Count[0]));
   CLKNAND2X2M U29 (.Y(n5), 
	.B(En), 
	.A(Samples[2]));
   MXI2X1M U30 (.Y(n24), 
	.S0(n21), 
	.B(n26), 
	.A(n6));
   NAND4X1M U31 (.Y(n21), 
	.D(n30), 
	.C(n29), 
	.B(n28), 
	.A(n27));
   NOR4BX1M U32 (.Y(n30), 
	.D(n32), 
	.C(n31), 
	.B(Edge_Count[5]), 
	.AN(n22));
   CLKXOR2X2M U33 (.Y(n32), 
	.B(Edge_Count[1]), 
	.A(Prescale[2]));
   CLKXOR2X2M U34 (.Y(n31), 
	.B(Edge_Count[0]), 
	.A(Prescale[1]));
   XNOR2X1M U35 (.Y(n29), 
	.B(Prescale[4]), 
	.A(Edge_Count[3]));
   CLKXOR2X2M U36 (.Y(n28), 
	.B(Prescale[5]), 
	.A(n19));
   CLKINVX1M U37 (.Y(n19), 
	.A(Edge_Count[4]));
   XNOR2X1M U38 (.Y(n27), 
	.B(Prescale[3]), 
	.A(Edge_Count[2]));
   CLKNAND2X2M U39 (.Y(n26), 
	.B(En), 
	.A(Samples[1]));
   MXI2X1M U40 (.Y(n23), 
	.S0(n22), 
	.B(n33), 
	.A(n6));
   NAND4X1M U41 (.Y(n22), 
	.D(n37), 
	.C(n36), 
	.B(n35), 
	.A(n34));
   NOR3X1M U42 (.Y(n37), 
	.C(n39), 
	.B(Edge_Count[5]), 
	.A(n38));
   CLKXOR2X2M U43 (.Y(n39), 
	.B(Edge_Count[0]), 
	.A(Middle_Sample_minus[0]));
   CLKXOR2X2M U44 (.Y(n38), 
	.B(Edge_Count[4]), 
	.A(Middle_Sample_minus[4]));
   XNOR2X1M U45 (.Y(n36), 
	.B(Middle_Sample_minus[2]), 
	.A(Edge_Count[2]));
   XNOR2X1M U46 (.Y(n35), 
	.B(Middle_Sample_minus[3]), 
	.A(Edge_Count[3]));
   CLKXOR2X2M U47 (.Y(n34), 
	.B(Middle_Sample_minus[1]), 
	.A(n18));
   CLKINVX1M U48 (.Y(n18), 
	.A(Edge_Count[1]));
   CLKNAND2X2M U49 (.Y(n33), 
	.B(En), 
	.A(Samples[0]));
   CLKNAND2X2M U50 (.Y(n6), 
	.B(En), 
	.A(RX_In));
   AOI21BX1M U51 (.Y(N25), 
	.B0N(En), 
	.A1(n41), 
	.A0(n40));
   OAI21X1M U52 (.Y(n41), 
	.B0(Samples[2]), 
	.A1(Samples[1]), 
	.A0(Samples[0]));
   CLKNAND2X2M U53 (.Y(n40), 
	.B(Samples[1]), 
	.A(Samples[0]));
endmodule

module Deserializer_Data_Width8_test_1 (
	CLK, 
	RST, 
	En, 
	Prescale, 
	S_In, 
	edge_count, 
	P_out, 
	Deser_Done, 
	test_si, 
	test_so, 
	test_se);
   input CLK;
   input RST;
   input En;
   input [5:0] Prescale;
   input S_In;
   input [5:0] edge_count;
   output [7:0] P_out;
   output Deser_Done;
   input test_si;
   output test_so;
   input test_se;

   // Internal wires
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire n15;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n17;
   wire n18;
   wire n19;
   wire n27;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n65;
   wire n66;
   wire [3:0] N;

   assign test_so = n20 ;

   SDFFRX1M \P_out_reg[5]  (.SI(n23), 
	.SE(n66), 
	.RN(RST), 
	.QN(n22), 
	.Q(P_out[5]), 
	.D(n41), 
	.CK(CLK));
   SDFFRX1M \P_out_reg[1]  (.SI(P_out[0]), 
	.SE(n66), 
	.RN(RST), 
	.QN(n26), 
	.Q(P_out[1]), 
	.D(n37), 
	.CK(CLK));
   SDFFRX1M \P_out_reg[4]  (.SI(n24), 
	.SE(n66), 
	.RN(RST), 
	.QN(n23), 
	.Q(P_out[4]), 
	.D(n40), 
	.CK(CLK));
   SDFFRQX2M \P_out_reg[0]  (.SI(n62), 
	.SE(n66), 
	.RN(RST), 
	.Q(P_out[0]), 
	.D(n36), 
	.CK(CLK));
   SDFFRX1M \P_out_reg[3]  (.SI(n25), 
	.SE(n66), 
	.RN(RST), 
	.QN(n24), 
	.Q(P_out[3]), 
	.D(n39), 
	.CK(CLK));
   SDFFRX1M \P_out_reg[2]  (.SI(n26), 
	.SE(n66), 
	.RN(RST), 
	.QN(n25), 
	.Q(P_out[2]), 
	.D(n38), 
	.CK(CLK));
   SDFFRX1M \P_out_reg[6]  (.SI(n22), 
	.SE(n66), 
	.RN(RST), 
	.QN(n21), 
	.Q(P_out[6]), 
	.D(n42), 
	.CK(CLK));
   SDFFRX1M \P_out_reg[7]  (.SI(n21), 
	.SE(n66), 
	.RN(RST), 
	.QN(n20), 
	.Q(P_out[7]), 
	.D(n43), 
	.CK(CLK));
   SDFFRQX2M \N_reg[0]  (.SI(test_si), 
	.SE(n66), 
	.RN(RST), 
	.Q(N[0]), 
	.D(n46), 
	.CK(CLK));
   SDFFRQX2M \N_reg[2]  (.SI(n60), 
	.SE(n66), 
	.RN(RST), 
	.Q(N[2]), 
	.D(n58), 
	.CK(CLK));
   SDFFRQX2M \N_reg[1]  (.SI(n59), 
	.SE(n66), 
	.RN(RST), 
	.Q(N[1]), 
	.D(n45), 
	.CK(CLK));
   SDFFRX1M \N_reg[3]  (.SI(n61), 
	.SE(n66), 
	.RN(RST), 
	.QN(n15), 
	.Q(n62), 
	.D(n44), 
	.CK(CLK));
   NOR2X2M U18 (.Y(n31), 
	.B(n28), 
	.A(n59));
   NAND2X2M U19 (.Y(n35), 
	.B(n28), 
	.A(En));
   INVX2M U20 (.Y(n57), 
	.A(n28));
   OAI21X2M U21 (.Y(n32), 
	.B0(n34), 
	.A1(n28), 
	.A0(N[1]));
   OAI22X1M U22 (.Y(n46), 
	.B1(n28), 
	.B0(N[0]), 
	.A1(n35), 
	.A0(n59));
   OAI22X1M U23 (.Y(n37), 
	.B1(n25), 
	.B0(n28), 
	.A1(n26), 
	.A0(n57));
   OAI22X1M U24 (.Y(n38), 
	.B1(n24), 
	.B0(n28), 
	.A1(n25), 
	.A0(n57));
   OAI22X1M U25 (.Y(n39), 
	.B1(n23), 
	.B0(n28), 
	.A1(n24), 
	.A0(n57));
   OAI22X1M U26 (.Y(n40), 
	.B1(n22), 
	.B0(n28), 
	.A1(n23), 
	.A0(n57));
   OAI22X1M U27 (.Y(n41), 
	.B1(n21), 
	.B0(n28), 
	.A1(n22), 
	.A0(n57));
   OAI22X1M U28 (.Y(n42), 
	.B1(n20), 
	.B0(n28), 
	.A1(n21), 
	.A0(n57));
   NAND2X2M U29 (.Y(n28), 
	.B(En), 
	.A(N10));
   OAI2BB2X1M U30 (.Y(n45), 
	.B1(n60), 
	.B0(n34), 
	.A1N(n31), 
	.A0N(n60));
   INVX2M U31 (.Y(n60), 
	.A(N[1]));
   OAI2BB2X1M U32 (.Y(n36), 
	.B1(n26), 
	.B0(n28), 
	.A1N(n28), 
	.A0N(P_out[0]));
   OR2X2M U33 (.Y(n17), 
	.B(Prescale[0]), 
	.A(Prescale[1]));
   OAI2BB2X1M U34 (.Y(n43), 
	.B1(n20), 
	.B0(n57), 
	.A1N(n57), 
	.A0N(S_In));
   OAI21X2M U35 (.Y(n44), 
	.B0(n30), 
	.A1(n15), 
	.A0(n29));
   NAND4X2M U36 (.Y(n30), 
	.D(n15), 
	.C(n31), 
	.B(N[1]), 
	.A(N[2]));
   AOI21X2M U37 (.Y(n29), 
	.B0(n32), 
	.A1(n61), 
	.A0(n57));
   OA21X2M U38 (.Y(n34), 
	.B0(n35), 
	.A1(n28), 
	.A0(N[0]));
   INVX2M U39 (.Y(n47), 
	.A(Prescale[3]));
   INVX2M U40 (.Y(n58), 
	.A(n33));
   AOI32X1M U41 (.Y(n33), 
	.B1(N[2]), 
	.B0(n32), 
	.A2(n31), 
	.A1(n61), 
	.A0(N[1]));
   NOR4X1M U42 (.Y(Deser_Done), 
	.D(n15), 
	.C(N[0]), 
	.B(N[1]), 
	.A(N[2]));
   INVX2M U43 (.Y(n59), 
	.A(N[0]));
   INVX2M U44 (.Y(n61), 
	.A(N[2]));
   CLKINVX1M U45 (.Y(N4), 
	.A(Prescale[0]));
   OAI2BB1X1M U46 (.Y(N5), 
	.B0(n17), 
	.A1N(Prescale[1]), 
	.A0N(Prescale[0]));
   NOR2X1M U47 (.Y(n18), 
	.B(Prescale[2]), 
	.A(n17));
   AO21XLM U48 (.Y(N6), 
	.B0(n18), 
	.A1(Prescale[2]), 
	.A0(n17));
   CLKNAND2X2M U49 (.Y(n19), 
	.B(n47), 
	.A(n18));
   OAI21X1M U50 (.Y(N7), 
	.B0(n19), 
	.A1(n47), 
	.A0(n18));
   XNOR2X1M U51 (.Y(N8), 
	.B(n19), 
	.A(Prescale[4]));
   NOR2X1M U52 (.Y(n27), 
	.B(n19), 
	.A(Prescale[4]));
   CLKXOR2X2M U53 (.Y(N9), 
	.B(n27), 
	.A(Prescale[5]));
   NOR2BX1M U54 (.Y(n48), 
	.B(N4), 
	.AN(edge_count[0]));
   OAI2B2X1M U55 (.Y(n52), 
	.B1(n48), 
	.B0(edge_count[1]), 
	.A1N(N5), 
	.A0(n48));
   NOR2BX1M U56 (.Y(n49), 
	.B(edge_count[0]), 
	.AN(N4));
   OAI2B2X1M U57 (.Y(n51), 
	.B1(n49), 
	.B0(N5), 
	.A1N(edge_count[1]), 
	.A0(n49));
   XNOR2X1M U58 (.Y(n50), 
	.B(edge_count[5]), 
	.A(N9));
   NAND3X1M U59 (.Y(n56), 
	.C(n50), 
	.B(n51), 
	.A(n52));
   CLKXOR2X2M U60 (.Y(n55), 
	.B(edge_count[4]), 
	.A(N8));
   CLKXOR2X2M U61 (.Y(n54), 
	.B(edge_count[2]), 
	.A(N6));
   CLKXOR2X2M U62 (.Y(n53), 
	.B(edge_count[3]), 
	.A(N7));
   NOR4X1M U63 (.Y(N10), 
	.D(n53), 
	.C(n54), 
	.B(n55), 
	.A(n56));
   INVXLM U64 (.Y(n65), 
	.A(test_se));
   CLKINVX2M U65 (.Y(n66), 
	.A(n65));
endmodule

module Edge_Bit_Counter_Data_Width8_test_1 (
	CLK, 
	RST, 
	En, 
	Prescale, 
	Bit_Count, 
	Edge_Count, 
	test_si, 
	test_se);
   input CLK;
   input RST;
   input En;
   input [5:0] Prescale;
   output [3:0] Bit_Count;
   output [5:0] Edge_Count;
   input test_si;
   input test_se;

   // Internal wires
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire \add_39/carry[5] ;
   wire \add_39/carry[4] ;
   wire \add_39/carry[3] ;
   wire \add_39/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;

   SDFFRQX2M \Bit_Count_reg[2]  (.SI(n38), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Bit_Count[2]), 
	.D(n29), 
	.CK(CLK));
   SDFFRQX2M \Bit_Count_reg[3]  (.SI(n39), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Bit_Count[3]), 
	.D(n28), 
	.CK(CLK));
   SDFFRQX2M \Bit_Count_reg[1]  (.SI(n37), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Bit_Count[1]), 
	.D(n30), 
	.CK(CLK));
   SDFFRQX2M \Bit_Count_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Bit_Count[0]), 
	.D(n31), 
	.CK(CLK));
   SDFFRQX2M \Edge_Count_reg[5]  (.SI(Edge_Count[4]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Edge_Count[5]), 
	.D(N32), 
	.CK(CLK));
   SDFFRQX2M \Edge_Count_reg[0]  (.SI(n40), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Edge_Count[0]), 
	.D(N27), 
	.CK(CLK));
   SDFFRQX2M \Edge_Count_reg[4]  (.SI(Edge_Count[3]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Edge_Count[4]), 
	.D(N31), 
	.CK(CLK));
   SDFFRQX2M \Edge_Count_reg[1]  (.SI(N15), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Edge_Count[1]), 
	.D(N28), 
	.CK(CLK));
   SDFFRQX2M \Edge_Count_reg[3]  (.SI(Edge_Count[2]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Edge_Count[3]), 
	.D(N30), 
	.CK(CLK));
   SDFFRQX2M \Edge_Count_reg[2]  (.SI(Edge_Count[1]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Edge_Count[2]), 
	.D(N29), 
	.CK(CLK));
   INVX2M U6 (.Y(n34), 
	.A(n27));
   INVX2M U7 (.Y(n35), 
	.A(En));
   NOR2X2M U15 (.Y(n27), 
	.B(N11), 
	.A(n35));
   AOI21X2M U16 (.Y(n26), 
	.B0(n27), 
	.A1(En), 
	.A0(n37));
   AND2X2M U17 (.Y(N28), 
	.B(n27), 
	.A(N16));
   AND2X2M U18 (.Y(N29), 
	.B(n27), 
	.A(N17));
   AND2X2M U19 (.Y(N30), 
	.B(n27), 
	.A(N18));
   AND2X2M U20 (.Y(N31), 
	.B(n27), 
	.A(N19));
   NOR3X2M U21 (.Y(n23), 
	.C(n39), 
	.B(n37), 
	.A(n38));
   OAI32X1M U22 (.Y(n31), 
	.B1(n34), 
	.B0(n37), 
	.A2(n27), 
	.A1(Bit_Count[0]), 
	.A0(n35));
   OAI32X1M U23 (.Y(n29), 
	.B1(n39), 
	.B0(n25), 
	.A2(n38), 
	.A1(Bit_Count[2]), 
	.A0(n24));
   OA21X2M U24 (.Y(n25), 
	.B0(n26), 
	.A1(Bit_Count[1]), 
	.A0(n35));
   OAI22X1M U25 (.Y(n28), 
	.B1(n35), 
	.B0(n22), 
	.A1(n34), 
	.A0(n40));
   AOI32X1M U26 (.Y(n22), 
	.B1(n36), 
	.B0(Bit_Count[3]), 
	.A2(N11), 
	.A1(n40), 
	.A0(n23));
   INVX2M U27 (.Y(n40), 
	.A(Bit_Count[3]));
   INVX2M U28 (.Y(n36), 
	.A(n23));
   NAND3X2M U29 (.Y(n24), 
	.C(En), 
	.B(n34), 
	.A(Bit_Count[0]));
   OAI22X1M U30 (.Y(n30), 
	.B1(n24), 
	.B0(Bit_Count[1]), 
	.A1(n38), 
	.A0(n26));
   OR2X2M U31 (.Y(n1), 
	.B(Prescale[0]), 
	.A(Prescale[1]));
   AND2X2M U32 (.Y(N32), 
	.B(n27), 
	.A(N20));
   AND2X2M U33 (.Y(N27), 
	.B(n27), 
	.A(N15));
   INVX2M U34 (.Y(n37), 
	.A(Bit_Count[0]));
   INVX2M U35 (.Y(n38), 
	.A(Bit_Count[1]));
   ADDHX1M U36 (.S(N17), 
	.CO(\add_39/carry[3] ), 
	.B(\add_39/carry[2] ), 
	.A(Edge_Count[2]));
   ADDHX1M U37 (.S(N18), 
	.CO(\add_39/carry[4] ), 
	.B(\add_39/carry[3] ), 
	.A(Edge_Count[3]));
   ADDHX1M U38 (.S(N16), 
	.CO(\add_39/carry[2] ), 
	.B(Edge_Count[0]), 
	.A(Edge_Count[1]));
   INVX2M U39 (.Y(n39), 
	.A(Bit_Count[2]));
   ADDHX1M U40 (.S(N19), 
	.CO(\add_39/carry[5] ), 
	.B(\add_39/carry[4] ), 
	.A(Edge_Count[4]));
   CLKINVX1M U41 (.Y(N4), 
	.A(Prescale[0]));
   OAI2BB1X1M U42 (.Y(N5), 
	.B0(n1), 
	.A1N(Prescale[1]), 
	.A0N(Prescale[0]));
   OR2X1M U43 (.Y(n2), 
	.B(Prescale[2]), 
	.A(n1));
   OAI2BB1X1M U44 (.Y(N6), 
	.B0(n2), 
	.A1N(Prescale[2]), 
	.A0N(n1));
   OR2X1M U45 (.Y(n3), 
	.B(Prescale[3]), 
	.A(n2));
   OAI2BB1X1M U46 (.Y(N7), 
	.B0(n3), 
	.A1N(Prescale[3]), 
	.A0N(n2));
   OR2X1M U47 (.Y(n4), 
	.B(Prescale[4]), 
	.A(n3));
   OAI2BB1X1M U48 (.Y(N8), 
	.B0(n4), 
	.A1N(Prescale[4]), 
	.A0N(n3));
   NOR2X1M U49 (.Y(N10), 
	.B(Prescale[5]), 
	.A(n4));
   AO21XLM U50 (.Y(N9), 
	.B0(N10), 
	.A1(Prescale[5]), 
	.A0(n4));
   CLKINVX1M U51 (.Y(N15), 
	.A(Edge_Count[0]));
   CLKXOR2X2M U52 (.Y(N20), 
	.B(Edge_Count[5]), 
	.A(\add_39/carry[5] ));
   NOR2BX1M U53 (.Y(n15), 
	.B(Edge_Count[0]), 
	.AN(N4));
   OAI2B2X1M U54 (.Y(n19), 
	.B1(n15), 
	.B0(N5), 
	.A1N(Edge_Count[1]), 
	.A0(n15));
   XNOR2X1M U55 (.Y(n18), 
	.B(Edge_Count[5]), 
	.A(N9));
   NOR2BX1M U56 (.Y(n16), 
	.B(N4), 
	.AN(Edge_Count[0]));
   OAI2B2X1M U57 (.Y(n17), 
	.B1(n16), 
	.B0(Edge_Count[1]), 
	.A1N(N5), 
	.A0(n16));
   NAND4BX1M U58 (.Y(n33), 
	.D(n17), 
	.C(n18), 
	.B(n19), 
	.AN(N10));
   CLKXOR2X2M U59 (.Y(n32), 
	.B(Edge_Count[4]), 
	.A(N8));
   CLKXOR2X2M U60 (.Y(n21), 
	.B(Edge_Count[2]), 
	.A(N6));
   CLKXOR2X2M U61 (.Y(n20), 
	.B(Edge_Count[3]), 
	.A(N7));
   NOR4X1M U62 (.Y(N11), 
	.D(n20), 
	.C(n21), 
	.B(n32), 
	.A(n33));
endmodule

module Parity_Check_Data_Width8_test_1 (
	CLK, 
	RST, 
	En, 
	Flags_Done, 
	PAR_TYP, 
	R_Data, 
	Deser_Done, 
	Parity_In, 
	par_err, 
	test_si, 
	test_se);
   input CLK;
   input RST;
   input En;
   input Flags_Done;
   input PAR_TYP;
   input [7:0] R_Data;
   input Deser_Done;
   input Parity_In;
   output par_err;
   input test_si;
   input test_se;

   // Internal wires
   wire Calc_parity;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n3;
   wire n4;

   SDFFRQX2M Calc_parity_reg (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Calc_parity), 
	.D(n14), 
	.CK(CLK));
   SDFFRQX2M par_err_reg (.SI(Calc_parity), 
	.SE(test_se), 
	.RN(RST), 
	.Q(par_err), 
	.D(n13), 
	.CK(CLK));
   NOR2X2M U5 (.Y(n7), 
	.B(En), 
	.A(Flags_Done));
   OAI31X1M U6 (.Y(n13), 
	.B0(n6), 
	.A2(n5), 
	.A1(Deser_Done), 
	.A0(n3));
   XNOR2X2M U7 (.Y(n5), 
	.B(Parity_In), 
	.A(Calc_parity));
   OAI21X2M U8 (.Y(n6), 
	.B0(par_err), 
	.A1(Deser_Done), 
	.A0(n7));
   INVX2M U9 (.Y(n3), 
	.A(En));
   XNOR2X2M U10 (.Y(n11), 
	.B(R_Data[2]), 
	.A(R_Data[3]));
   XOR3XLM U11 (.Y(n9), 
	.C(n12), 
	.B(R_Data[4]), 
	.A(R_Data[5]));
   CLKXOR2X2M U12 (.Y(n12), 
	.B(R_Data[6]), 
	.A(R_Data[7]));
   OAI2BB2X1M U13 (.Y(n14), 
	.B1(n4), 
	.B0(n8), 
	.A1N(Calc_parity), 
	.A0N(n4));
   INVX2M U14 (.Y(n4), 
	.A(Deser_Done));
   XOR3XLM U15 (.Y(n8), 
	.C(n10), 
	.B(PAR_TYP), 
	.A(n9));
   XOR3XLM U16 (.Y(n10), 
	.C(n11), 
	.B(R_Data[0]), 
	.A(R_Data[1]));
endmodule

module Start_Check_test_1 (
	CLK, 
	RST, 
	En, 
	Start_bit, 
	Str_err, 
	test_si, 
	test_se);
   input CLK;
   input RST;
   input En;
   input Start_bit;
   output Str_err;
   input test_si;
   input test_se;

   // Internal wires
   wire N4;

   SDFFRQX2M Str_err_reg (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Str_err), 
	.D(N4), 
	.CK(CLK));
   AND2X2M U4 (.Y(N4), 
	.B(En), 
	.A(Start_bit));
endmodule

module Stop_Check_test_1 (
	CLK, 
	RST, 
	En, 
	Flags_Done, 
	Stop_bit, 
	Stp_err, 
	test_si, 
	test_so, 
	test_se);
   input CLK;
   input RST;
   input En;
   input Flags_Done;
   input Stop_bit;
   output Stp_err;
   input test_si;
   output test_so;
   input test_se;

   // Internal wires
   wire n2;
   wire n4;
   wire n3;

   assign test_so = n2 ;

   SDFFRX1M Stp_err_reg (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.QN(n2), 
	.Q(Stp_err), 
	.D(n4), 
	.CK(CLK));
   OAI32X1M U4 (.Y(n4), 
	.B1(n3), 
	.B0(Stop_bit), 
	.A2(En), 
	.A1(Flags_Done), 
	.A0(n2));
   INVX2M U5 (.Y(n3), 
	.A(En));
endmodule

module RX_FSM_Data_Width8_test_1 (
	CLK, 
	RST, 
	PAR_EN, 
	Prescale, 
	RX_In, 
	Bit_Count, 
	edge_count, 
	Par_err, 
	Start_err, 
	Stop_err, 
	edge_bit_en, 
	data_samp_en, 
	Deser_en, 
	Par_chk_en, 
	Str_chk_en, 
	Stp_chk_en, 
	Flags_Done, 
	Parity_Error, 
	Stop_Error, 
	Data_Valid, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN5_M_Domain2_SYNC_RST, 
	RX_CLK_M__L3_N1);
   input CLK;
   input RST;
   input PAR_EN;
   input [5:0] Prescale;
   input RX_In;
   input [3:0] Bit_Count;
   input [5:0] edge_count;
   input Par_err;
   input Start_err;
   input Stop_err;
   output edge_bit_en;
   output data_samp_en;
   output Deser_en;
   output Par_chk_en;
   output Str_chk_en;
   output Stp_chk_en;
   output Flags_Done;
   output Parity_Error;
   output Stop_Error;
   output Data_Valid;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN5_M_Domain2_SYNC_RST;
   input RX_CLK_M__L3_N1;

   // Internal wires
   wire Parity_Error_c;
   wire Stop_Error_c;
   wire Data_Valid_c;
   wire \add_78/carry[4] ;
   wire \add_78/carry[3] ;
   wire \sub_77/carry[5] ;
   wire \sub_77/carry[4] ;
   wire \sub_77/carry[3] ;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire [5:0] Final_edge;
   wire [5:0] Flags_edge;
   wire [5:0] Check_edge;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign Flags_edge[0] = Prescale[0] ;
   assign Check_edge[0] = Prescale[1] ;
   assign test_so = current_state[2] ;

   SDFFRQX2M \current_state_reg[2]  (.SI(current_state[1]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(current_state[2]), 
	.D(next_state[2]), 
	.CK(RX_CLK_M__L3_N1));
   SDFFRQX2M \current_state_reg[0]  (.SI(Stop_Error), 
	.SE(test_se), 
	.RN(RST), 
	.Q(current_state[0]), 
	.D(next_state[0]), 
	.CK(RX_CLK_M__L3_N1));
   SDFFRQX2M \current_state_reg[1]  (.SI(current_state[0]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(current_state[1]), 
	.D(next_state[1]), 
	.CK(RX_CLK_M__L3_N1));
   SDFFRQX4M Stop_Error_reg (.SI(Parity_Error), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Stop_Error), 
	.D(Stop_Error_c), 
	.CK(CLK));
   SDFFRQX4M Parity_Error_reg (.SI(Data_Valid), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Parity_Error), 
	.D(Parity_Error_c), 
	.CK(CLK));
   SDFFRQX2M Data_Valid_reg (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Data_Valid), 
	.D(Data_Valid_c), 
	.CK(RX_CLK_M__L3_N1));
   INVX2M U7 (.Y(Check_edge[1]), 
	.A(Prescale[2]));
   OR2X2M U8 (.Y(n2), 
	.B(Flags_edge[0]), 
	.A(Check_edge[0]));
   INVX2M U9 (.Y(n6), 
	.A(Prescale[3]));
   INVX2M U10 (.Y(Flags_edge[1]), 
	.A(Check_edge[0]));
   XNOR2X1M U14 (.Y(Flags_edge[5]), 
	.B(\sub_77/carry[5] ), 
	.A(Prescale[5]));
   OR2X1M U15 (.Y(\sub_77/carry[5] ), 
	.B(\sub_77/carry[4] ), 
	.A(Prescale[4]));
   XNOR2X1M U16 (.Y(Flags_edge[4]), 
	.B(Prescale[4]), 
	.A(\sub_77/carry[4] ));
   OR2X1M U17 (.Y(\sub_77/carry[4] ), 
	.B(\sub_77/carry[3] ), 
	.A(Prescale[3]));
   XNOR2X1M U18 (.Y(Flags_edge[3]), 
	.B(Prescale[3]), 
	.A(\sub_77/carry[3] ));
   OR2X1M U19 (.Y(\sub_77/carry[3] ), 
	.B(Check_edge[0]), 
	.A(Prescale[2]));
   XNOR2X1M U20 (.Y(Flags_edge[2]), 
	.B(Prescale[2]), 
	.A(Check_edge[0]));
   AND2X1M U21 (.Y(Check_edge[5]), 
	.B(Prescale[5]), 
	.A(\add_78/carry[4] ));
   CLKXOR2X2M U22 (.Y(Check_edge[4]), 
	.B(\add_78/carry[4] ), 
	.A(Prescale[5]));
   AND2X1M U23 (.Y(\add_78/carry[4] ), 
	.B(Prescale[4]), 
	.A(\add_78/carry[3] ));
   CLKXOR2X2M U24 (.Y(Check_edge[3]), 
	.B(\add_78/carry[3] ), 
	.A(Prescale[4]));
   AND2X1M U25 (.Y(\add_78/carry[3] ), 
	.B(Prescale[3]), 
	.A(Prescale[2]));
   CLKXOR2X2M U26 (.Y(Check_edge[2]), 
	.B(Prescale[2]), 
	.A(Prescale[3]));
   CLKINVX1M U27 (.Y(Final_edge[0]), 
	.A(Flags_edge[0]));
   OAI2BB1X1M U28 (.Y(Final_edge[1]), 
	.B0(n2), 
	.A1N(Check_edge[0]), 
	.A0N(Flags_edge[0]));
   NOR2X1M U29 (.Y(n3), 
	.B(Prescale[2]), 
	.A(n2));
   AO21XLM U30 (.Y(Final_edge[2]), 
	.B0(n3), 
	.A1(Prescale[2]), 
	.A0(n2));
   CLKNAND2X2M U31 (.Y(n4), 
	.B(n6), 
	.A(n3));
   OAI21X1M U32 (.Y(Final_edge[3]), 
	.B0(n4), 
	.A1(n6), 
	.A0(n3));
   XNOR2X1M U33 (.Y(Final_edge[4]), 
	.B(n4), 
	.A(Prescale[4]));
   NOR2X1M U34 (.Y(n5), 
	.B(n4), 
	.A(Prescale[4]));
   CLKXOR2X2M U35 (.Y(Final_edge[5]), 
	.B(n5), 
	.A(Prescale[5]));
   OAI32X1M U36 (.Y(next_state[2]), 
	.B1(n11), 
	.B0(n10), 
	.A2(n9), 
	.A1(n8), 
	.A0(n7));
   MXI2X1M U37 (.Y(n7), 
	.S0(Bit_Count[0]), 
	.B(n13), 
	.A(n12));
   NOR2X1M U38 (.Y(n12), 
	.B(n14), 
	.A(PAR_EN));
   OAI21X1M U39 (.Y(next_state[1]), 
	.B0(n22), 
	.A1(n15), 
	.A0(current_state[2]));
   AOI32X1M U40 (.Y(n22), 
	.B1(n26), 
	.B0(n13), 
	.A2(n25), 
	.A1(n24), 
	.A0(n23));
   NAND4X1M U41 (.Y(n26), 
	.D(n30), 
	.C(n29), 
	.B(n28), 
	.A(n27));
   NOR4X1M U42 (.Y(n30), 
	.D(n34), 
	.C(n33), 
	.B(n32), 
	.A(n31));
   CLKXOR2X2M U43 (.Y(n34), 
	.B(Flags_edge[5]), 
	.A(edge_count[5]));
   CLKXOR2X2M U44 (.Y(n33), 
	.B(Flags_edge[4]), 
	.A(edge_count[4]));
   CLKXOR2X2M U45 (.Y(n32), 
	.B(Flags_edge[3]), 
	.A(edge_count[3]));
   CLKXOR2X2M U46 (.Y(n31), 
	.B(Flags_edge[2]), 
	.A(edge_count[2]));
   NOR3X1M U47 (.Y(n29), 
	.C(n35), 
	.B(Bit_Count[2]), 
	.A(n9));
   XNOR2X1M U48 (.Y(n35), 
	.B(Bit_Count[0]), 
	.A(Bit_Count[1]));
   CLKINVX1M U49 (.Y(n9), 
	.A(Bit_Count[3]));
   CLKXOR2X2M U50 (.Y(n28), 
	.B(Flags_edge[0]), 
	.A(n36));
   CLKINVX1M U51 (.Y(n36), 
	.A(edge_count[0]));
   CLKXOR2X2M U52 (.Y(n27), 
	.B(Flags_edge[1]), 
	.A(n37));
   CLKINVX1M U53 (.Y(n37), 
	.A(edge_count[1]));
   NOR3X1M U54 (.Y(n25), 
	.C(Bit_Count[3]), 
	.B(Start_err), 
	.A(Bit_Count[0]));
   CLKINVX1M U55 (.Y(n23), 
	.A(n8));
   OAI211X1M U56 (.Y(next_state[0]), 
	.C0(n39), 
	.B0(n38), 
	.A1(n14), 
	.A0(Bit_Count[3]));
   OR3X1M U57 (.Y(n39), 
	.C(current_state[0]), 
	.B(current_state[1]), 
	.A(RX_In));
   OAI31X1M U58 (.Y(n38), 
	.B0(n24), 
	.A2(n8), 
	.A1(Bit_Count[0]), 
	.A0(n40));
   CLKNAND2X2M U59 (.Y(n8), 
	.B(n42), 
	.A(n41));
   NOR4X1M U60 (.Y(n42), 
	.D(n44), 
	.C(n43), 
	.B(Bit_Count[1]), 
	.A(Bit_Count[2]));
   CLKXOR2X2M U61 (.Y(n44), 
	.B(Final_edge[0]), 
	.A(edge_count[0]));
   CLKXOR2X2M U62 (.Y(n43), 
	.B(Final_edge[4]), 
	.A(edge_count[4]));
   NOR4X1M U63 (.Y(n41), 
	.D(n48), 
	.C(n47), 
	.B(n46), 
	.A(n45));
   CLKXOR2X2M U64 (.Y(n48), 
	.B(Final_edge[3]), 
	.A(edge_count[3]));
   CLKXOR2X2M U65 (.Y(n47), 
	.B(Final_edge[2]), 
	.A(edge_count[2]));
   CLKXOR2X2M U66 (.Y(n46), 
	.B(Final_edge[5]), 
	.A(edge_count[5]));
   CLKXOR2X2M U67 (.Y(n45), 
	.B(Final_edge[1]), 
	.A(edge_count[1]));
   MXI2X1M U68 (.Y(n40), 
	.S0(Bit_Count[3]), 
	.B(current_state[1]), 
	.A(Start_err));
   CLKNAND2X2M U69 (.Y(edge_bit_en), 
	.B(n10), 
	.A(n49));
   NOR3X1M U70 (.Y(Str_chk_en), 
	.C(n49), 
	.B(current_state[1]), 
	.A(n50));
   NOR3X1M U71 (.Y(Stp_chk_en), 
	.C(n11), 
	.B(n10), 
	.A(n50));
   AND2X1M U72 (.Y(Stop_Error_c), 
	.B(Stop_err), 
	.A(Flags_Done));
   AND2X1M U73 (.Y(Parity_Error_c), 
	.B(Par_err), 
	.A(Flags_Done));
   NOR3X1M U74 (.Y(Par_chk_en), 
	.C(n10), 
	.B(current_state[2]), 
	.A(n50));
   CLKINVX1M U75 (.Y(n10), 
	.A(n13));
   NOR2X1M U76 (.Y(n13), 
	.B(current_state[0]), 
	.A(n15));
   CLKINVX1M U77 (.Y(n15), 
	.A(current_state[1]));
   NAND4X1M U78 (.Y(n50), 
	.D(n54), 
	.C(n53), 
	.B(n52), 
	.A(n51));
   NOR3X1M U79 (.Y(n54), 
	.C(n57), 
	.B(n56), 
	.A(n55));
   CLKXOR2X2M U80 (.Y(n57), 
	.B(Check_edge[4]), 
	.A(edge_count[4]));
   CLKXOR2X2M U81 (.Y(n56), 
	.B(Check_edge[1]), 
	.A(edge_count[1]));
   CLKXOR2X2M U82 (.Y(n55), 
	.B(Check_edge[0]), 
	.A(edge_count[0]));
   XNOR2X1M U83 (.Y(n53), 
	.B(Check_edge[2]), 
	.A(edge_count[2]));
   XNOR2X1M U84 (.Y(n52), 
	.B(Check_edge[3]), 
	.A(edge_count[3]));
   XNOR2X1M U85 (.Y(n51), 
	.B(Check_edge[5]), 
	.A(edge_count[5]));
   CLKINVX1M U86 (.Y(Deser_en), 
	.A(n14));
   CLKNAND2X2M U87 (.Y(n14), 
	.B(n24), 
	.A(current_state[1]));
   CLKINVX1M U88 (.Y(n24), 
	.A(n49));
   CLKNAND2X2M U89 (.Y(n49), 
	.B(n11), 
	.A(current_state[0]));
   NOR3BX1M U90 (.Y(Data_Valid_c), 
	.C(Par_err), 
	.B(Stop_err), 
	.AN(Flags_Done));
   NOR3X1M U91 (.Y(Flags_Done), 
	.C(n11), 
	.B(current_state[1]), 
	.A(current_state[0]));
   CLKINVX1M U92 (.Y(n11), 
	.A(current_state[2]));
endmodule

module UART_RX_TOP_Data_Width8_test_1 (
	CLK, 
	RST, 
	PAR_EN, 
	Prescale, 
	PAR_TYP, 
	RX_IN, 
	Paerity_Error, 
	Stop_Error, 
	Data_Valid, 
	P_DATA, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN5_M_Domain2_SYNC_RST, 
	RX_CLK_M__L3_N1);
   input CLK;
   input RST;
   input PAR_EN;
   input [5:0] Prescale;
   input PAR_TYP;
   input RX_IN;
   output Paerity_Error;
   output Stop_Error;
   output Data_Valid;
   output [7:0] P_DATA;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN5_M_Domain2_SYNC_RST;
   input RX_CLK_M__L3_N1;

   // Internal wires
   wire FE_PT0_;
   wire FE_UNCONNECTED_0;
   wire sampled_bit;
   wire deser_en;
   wire Deser_Done;
   wire edge_bit_en;
   wire Par_chk_en;
   wire Flags_Done;
   wire par_err;
   wire strt_chk_en;
   wire strt_glitch;
   wire stp_chk_en;
   wire stp_err;
   wire n4;
   wire n5;
   wire n6;
   wire [5:0] edge_cnt;
   wire [3:0] bit_cnt;

   Data_Sampling_test_1 U1 (.CLK(CLK), 
	.RST(RST), 
	.En(edge_bit_en), 
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }), 
	.RX_In(RX_IN), 
	.Edge_Count({ edge_cnt[5],
		edge_cnt[4],
		edge_cnt[3],
		edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }), 
	.Sampeld_Bit(sampled_bit), 
	.test_si(test_si), 
	.test_so(n6), 
	.test_se(test_se), 
	.RX_CLK_M__L3_N1(RX_CLK_M__L3_N1));
   Deserializer_Data_Width8_test_1 U2 (.CLK(CLK), 
	.RST(RST), 
	.En(deser_en), 
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }), 
	.S_In(sampled_bit), 
	.edge_count({ edge_cnt[5],
		edge_cnt[4],
		edge_cnt[3],
		edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }), 
	.P_out({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }), 
	.Deser_Done(Deser_Done), 
	.test_si(n6), 
	.test_so(n5), 
	.test_se(test_se));
   Edge_Bit_Counter_Data_Width8_test_1 U3 (.CLK(RX_CLK_M__L3_N1), 
	.RST(FE_OFN5_M_Domain2_SYNC_RST), 
	.En(edge_bit_en), 
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }), 
	.Bit_Count({ bit_cnt[3],
		bit_cnt[2],
		bit_cnt[1],
		bit_cnt[0] }), 
	.Edge_Count({ edge_cnt[5],
		edge_cnt[4],
		edge_cnt[3],
		edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }), 
	.test_si(n5), 
	.test_se(test_se));
   Parity_Check_Data_Width8_test_1 U4 (.CLK(CLK), 
	.RST(RST), 
	.En(Par_chk_en), 
	.Flags_Done(Flags_Done), 
	.PAR_TYP(PAR_TYP), 
	.R_Data({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }), 
	.Deser_Done(Deser_Done), 
	.Parity_In(sampled_bit), 
	.par_err(par_err), 
	.test_si(edge_cnt[5]), 
	.test_se(test_se));
   Start_Check_test_1 U5 (.CLK(RX_CLK_M__L3_N1), 
	.RST(FE_OFN5_M_Domain2_SYNC_RST), 
	.En(strt_chk_en), 
	.Start_bit(sampled_bit), 
	.Str_err(strt_glitch), 
	.test_si(par_err), 
	.test_se(test_se));
   Stop_Check_test_1 U6 (.CLK(RX_CLK_M__L3_N1), 
	.RST(FE_OFN5_M_Domain2_SYNC_RST), 
	.En(stp_chk_en), 
	.Flags_Done(Flags_Done), 
	.Stop_bit(sampled_bit), 
	.Stp_err(stp_err), 
	.test_si(strt_glitch), 
	.test_so(n4), 
	.test_se(test_se));
   RX_FSM_Data_Width8_test_1 U7 (.CLK(CLK), 
	.RST(RST), 
	.PAR_EN(PAR_EN), 
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }), 
	.RX_In(RX_IN), 
	.Bit_Count({ bit_cnt[3],
		bit_cnt[2],
		bit_cnt[1],
		bit_cnt[0] }), 
	.edge_count({ edge_cnt[5],
		edge_cnt[4],
		edge_cnt[3],
		edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }), 
	.Par_err(par_err), 
	.Start_err(strt_glitch), 
	.Stop_err(stp_err), 
	.edge_bit_en(edge_bit_en), 
	.data_samp_en(FE_PT0_), 
	.Deser_en(deser_en), 
	.Par_chk_en(Par_chk_en), 
	.Str_chk_en(strt_chk_en), 
	.Stp_chk_en(stp_chk_en), 
	.Flags_Done(Flags_Done), 
	.Parity_Error(Paerity_Error), 
	.Stop_Error(Stop_Error), 
	.Data_Valid(Data_Valid), 
	.test_si(n4), 
	.test_so(test_so), 
	.test_se(test_se), 
	.FE_OFN5_M_Domain2_SYNC_RST(FE_OFN5_M_Domain2_SYNC_RST), 
	.RX_CLK_M__L3_N1(RX_CLK_M__L3_N1));
endmodule

module MUX_4x1_test_1 (
	CLK, 
	RST, 
	mux_sel, 
	input_1, 
	input_2, 
	input_3, 
	input_4, 
	OUT, 
	test_si, 
	test_se);
   input CLK;
   input RST;
   input [1:0] mux_sel;
   input input_1;
   input input_2;
   input input_3;
   input input_4;
   output OUT;
   input test_si;
   input test_se;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire mux_out;
   wire n3;
   wire n4;
   wire n5;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   TIELOM LTIE_LTIELO (.Y(LTIE_LTIELO_NET));
   OAI2B2X1M U5 (.Y(mux_out), 
	.B1(n4), 
	.B0(mux_sel[1]), 
	.A1N(mux_sel[1]), 
	.A0(n3));
   AOI22X1M U6 (.Y(n4), 
	.B1(HTIE_LTIEHI_NET), 
	.B0(mux_sel[0]), 
	.A1(n5), 
	.A0(LTIE_LTIELO_NET));
   AOI22X1M U7 (.Y(n3), 
	.B1(mux_sel[0]), 
	.B0(input_4), 
	.A1(n5), 
	.A0(input_3));
   INVX2M U8 (.Y(n5), 
	.A(mux_sel[0]));
   SDFFSQX4M OUT_reg (.SN(RST), 
	.SI(test_si), 
	.SE(test_se), 
	.Q(OUT), 
	.D(mux_out), 
	.CK(CLK));
endmodule

module Parity_Calc_test_1 (
	CLK, 
	RST, 
	In_Data, 
	Data_Valid, 
	Basy_signal, 
	Parity_Calc_En, 
	PAR_TYP, 
	par_bit, 
	test_si, 
	test_se, 
	TX_CLK_M__L3_N1, 
	TX_CLK_M__L3_N2);
   input CLK;
   input RST;
   input [7:0] In_Data;
   input Data_Valid;
   input Basy_signal;
   input Parity_Calc_En;
   input PAR_TYP;
   output par_bit;
   input test_si;
   input test_se;
   input TX_CLK_M__L3_N1;
   input TX_CLK_M__L3_N2;

   // Internal wires
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire [7:0] DATA_V;

   SDFFRQX2M par_bit_reg (.SI(DATA_V[7]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(par_bit), 
	.D(n17), 
	.CK(CLK));
   SDFFRQX2M \DATA_V_reg[5]  (.SI(DATA_V[4]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(DATA_V[5]), 
	.D(n23), 
	.CK(TX_CLK_M__L3_N2));
   SDFFRQX2M \DATA_V_reg[1]  (.SI(DATA_V[0]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(DATA_V[1]), 
	.D(n19), 
	.CK(TX_CLK_M__L3_N1));
   SDFFRQX2M \DATA_V_reg[4]  (.SI(DATA_V[3]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(DATA_V[4]), 
	.D(n22), 
	.CK(TX_CLK_M__L3_N2));
   SDFFRQX2M \DATA_V_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.Q(DATA_V[0]), 
	.D(n18), 
	.CK(TX_CLK_M__L3_N1));
   SDFFRQX2M \DATA_V_reg[2]  (.SI(DATA_V[1]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(DATA_V[2]), 
	.D(n20), 
	.CK(TX_CLK_M__L3_N2));
   SDFFRQX2M \DATA_V_reg[3]  (.SI(DATA_V[2]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(DATA_V[3]), 
	.D(n21), 
	.CK(TX_CLK_M__L3_N2));
   SDFFRQX2M \DATA_V_reg[6]  (.SI(DATA_V[5]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(DATA_V[6]), 
	.D(n24), 
	.CK(TX_CLK_M__L3_N2));
   SDFFRQX2M \DATA_V_reg[7]  (.SI(DATA_V[6]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(DATA_V[7]), 
	.D(n25), 
	.CK(TX_CLK_M__L3_N1));
   NOR2BX2M U12 (.Y(n12), 
	.B(Basy_signal), 
	.AN(Data_Valid));
   XNOR2X2M U13 (.Y(n15), 
	.B(DATA_V[3]), 
	.A(DATA_V[2]));
   XOR3XLM U14 (.Y(n13), 
	.C(n16), 
	.B(DATA_V[4]), 
	.A(DATA_V[5]));
   CLKXOR2X2M U15 (.Y(n16), 
	.B(DATA_V[6]), 
	.A(DATA_V[7]));
   OAI2BB2X1M U16 (.Y(n17), 
	.B1(n11), 
	.B0(n10), 
	.A1N(n11), 
	.A0N(par_bit));
   XOR3XLM U17 (.Y(n10), 
	.C(n14), 
	.B(PAR_TYP), 
	.A(n13));
   NAND2BX2M U18 (.Y(n11), 
	.B(Parity_Calc_En), 
	.AN(n12));
   XOR3XLM U19 (.Y(n14), 
	.C(n15), 
	.B(DATA_V[0]), 
	.A(DATA_V[1]));
   AO2B2X2M U20 (.Y(n18), 
	.B1(n12), 
	.B0(In_Data[0]), 
	.A1N(n12), 
	.A0(DATA_V[0]));
   AO2B2X2M U21 (.Y(n19), 
	.B1(n12), 
	.B0(In_Data[1]), 
	.A1N(n12), 
	.A0(DATA_V[1]));
   AO2B2X2M U22 (.Y(n20), 
	.B1(n12), 
	.B0(In_Data[2]), 
	.A1N(n12), 
	.A0(DATA_V[2]));
   AO2B2X2M U23 (.Y(n21), 
	.B1(n12), 
	.B0(In_Data[3]), 
	.A1N(n12), 
	.A0(DATA_V[3]));
   AO2B2X2M U24 (.Y(n22), 
	.B1(n12), 
	.B0(In_Data[4]), 
	.A1N(n12), 
	.A0(DATA_V[4]));
   AO2B2X2M U25 (.Y(n23), 
	.B1(n12), 
	.B0(In_Data[5]), 
	.A1N(n12), 
	.A0(DATA_V[5]));
   AO2B2X2M U26 (.Y(n24), 
	.B1(n12), 
	.B0(In_Data[6]), 
	.A1N(n12), 
	.A0(DATA_V[6]));
   AO2B2X2M U27 (.Y(n25), 
	.B1(n12), 
	.B0(In_Data[7]), 
	.A1N(n12), 
	.A0(DATA_V[7]));
endmodule

module Serializer_1byte_test_1 (
	In_Data, 
	Data_Valid, 
	Basy_signal, 
	CLK, 
	RST, 
	ser_en, 
	ser_done, 
	Out_Data, 
	test_si, 
	test_se, 
	FE_OFN5_M_Domain2_SYNC_RST, 
	TX_CLK_M__L3_N1, 
	TX_CLK_M__L3_N2, 
	TX_CLK_M__L3_N3);
   input [7:0] In_Data;
   input Data_Valid;
   input Basy_signal;
   input CLK;
   input RST;
   input ser_en;
   output ser_done;
   output Out_Data;
   input test_si;
   input test_se;
   input FE_OFN5_M_Domain2_SYNC_RST;
   input TX_CLK_M__L3_N1;
   input TX_CLK_M__L3_N2;
   input TX_CLK_M__L3_N3;

   // Internal wires
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n48;
   wire [7:1] S_R_Data;
   wire [3:0] counter;

   SDFFRQX2M \S_R_Data_reg[6]  (.SI(S_R_Data[5]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(S_R_Data[6]), 
	.D(n38), 
	.CK(TX_CLK_M__L3_N1));
   SDFFRQX2M \S_R_Data_reg[5]  (.SI(S_R_Data[4]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(S_R_Data[5]), 
	.D(n39), 
	.CK(TX_CLK_M__L3_N1));
   SDFFRQX2M \S_R_Data_reg[4]  (.SI(S_R_Data[3]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(S_R_Data[4]), 
	.D(n40), 
	.CK(TX_CLK_M__L3_N3));
   SDFFRQX2M \S_R_Data_reg[3]  (.SI(S_R_Data[2]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(S_R_Data[3]), 
	.D(n41), 
	.CK(TX_CLK_M__L3_N2));
   SDFFRQX2M \S_R_Data_reg[2]  (.SI(S_R_Data[1]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(S_R_Data[2]), 
	.D(n42), 
	.CK(TX_CLK_M__L3_N1));
   SDFFRQX2M \S_R_Data_reg[1]  (.SI(Out_Data), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(S_R_Data[1]), 
	.D(n43), 
	.CK(TX_CLK_M__L3_N1));
   SDFFRQX2M \S_R_Data_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Out_Data), 
	.D(n36), 
	.CK(TX_CLK_M__L3_N1));
   SDFFRQX2M \S_R_Data_reg[7]  (.SI(S_R_Data[6]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(S_R_Data[7]), 
	.D(n37), 
	.CK(TX_CLK_M__L3_N1));
   SDFFRQX2M \counter_reg[3]  (.SI(counter[2]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(counter[3]), 
	.D(n46), 
	.CK(CLK));
   SDFFRQX2M \counter_reg[1]  (.SI(n18), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(counter[1]), 
	.D(n45), 
	.CK(TX_CLK_M__L3_N1));
   SDFFRQX2M \counter_reg[0]  (.SI(S_R_Data[7]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(counter[0]), 
	.D(n47), 
	.CK(TX_CLK_M__L3_N1));
   SDFFRQX2M \counter_reg[2]  (.SI(n48), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(counter[2]), 
	.D(n44), 
	.CK(CLK));
   SDFFRQX2M ser_done_reg (.SI(counter[3]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(ser_done), 
	.D(n15), 
	.CK(CLK));
   NOR2X2M U16 (.Y(n19), 
	.B(n16), 
	.A(n17));
   OAI21X2M U18 (.Y(n31), 
	.B0(n32), 
	.A1(n48), 
	.A0(n33));
   OAI21X2M U19 (.Y(n45), 
	.B0(n30), 
	.A1(n48), 
	.A0(n32));
   NAND3X2M U20 (.Y(n30), 
	.C(n17), 
	.B(n48), 
	.A(n18));
   INVX2M U21 (.Y(n17), 
	.A(n33));
   INVX2M U22 (.Y(n16), 
	.A(n35));
   NAND2X2M U23 (.Y(n29), 
	.B(n18), 
	.A(n28));
   AOI21X2M U24 (.Y(n32), 
	.B0(n19), 
	.A1(counter[0]), 
	.A0(n17));
   NAND2X2M U25 (.Y(n33), 
	.B(n35), 
	.A(ser_en));
   OAI211X2M U26 (.Y(n46), 
	.C0(n35), 
	.B0(n34), 
	.A1(n29), 
	.A0(n33));
   OAI21X2M U27 (.Y(n34), 
	.B0(counter[3]), 
	.A1(n31), 
	.A0(counter[2]));
   NAND2BX2M U28 (.Y(n35), 
	.B(Data_Valid), 
	.AN(Basy_signal));
   OAI2BB2X1M U29 (.Y(n44), 
	.B1(n30), 
	.B0(counter[2]), 
	.A1N(counter[2]), 
	.A0N(n31));
   OAI2BB2X1M U30 (.Y(n47), 
	.B1(n33), 
	.B0(counter[0]), 
	.A1N(counter[0]), 
	.A0N(n19));
   INVX2M U31 (.Y(n15), 
	.A(n27));
   AOI32X1M U32 (.Y(n27), 
	.B1(ser_done), 
	.B0(n19), 
	.A2(n17), 
	.A1(n29), 
	.A0(n28));
   OAI2BB1X2M U33 (.Y(n36), 
	.B0(n20), 
	.A1N(n19), 
	.A0N(Out_Data));
   AOI22X1M U34 (.Y(n20), 
	.B1(n17), 
	.B0(S_R_Data[1]), 
	.A1(n16), 
	.A0(In_Data[0]));
   OAI2BB1X2M U35 (.Y(n43), 
	.B0(n26), 
	.A1N(n19), 
	.A0N(S_R_Data[1]));
   AOI22X1M U36 (.Y(n26), 
	.B1(n17), 
	.B0(S_R_Data[2]), 
	.A1(n16), 
	.A0(In_Data[1]));
   OAI2BB1X2M U37 (.Y(n42), 
	.B0(n25), 
	.A1N(S_R_Data[2]), 
	.A0N(n19));
   AOI22X1M U38 (.Y(n25), 
	.B1(n17), 
	.B0(S_R_Data[3]), 
	.A1(n16), 
	.A0(In_Data[2]));
   OAI2BB1X2M U39 (.Y(n41), 
	.B0(n24), 
	.A1N(S_R_Data[3]), 
	.A0N(n19));
   AOI22X1M U40 (.Y(n24), 
	.B1(n17), 
	.B0(S_R_Data[4]), 
	.A1(n16), 
	.A0(In_Data[3]));
   OAI2BB1X2M U41 (.Y(n40), 
	.B0(n23), 
	.A1N(S_R_Data[4]), 
	.A0N(n19));
   AOI22X1M U42 (.Y(n23), 
	.B1(n17), 
	.B0(S_R_Data[5]), 
	.A1(n16), 
	.A0(In_Data[4]));
   OAI2BB1X2M U43 (.Y(n39), 
	.B0(n22), 
	.A1N(S_R_Data[5]), 
	.A0N(n19));
   AOI22X1M U44 (.Y(n22), 
	.B1(n17), 
	.B0(S_R_Data[6]), 
	.A1(n16), 
	.A0(In_Data[5]));
   OAI2BB1X2M U45 (.Y(n38), 
	.B0(n21), 
	.A1N(S_R_Data[6]), 
	.A0N(n19));
   AOI22X1M U46 (.Y(n21), 
	.B1(n17), 
	.B0(S_R_Data[7]), 
	.A1(n16), 
	.A0(In_Data[6]));
   AO22X1M U47 (.Y(n37), 
	.B1(n16), 
	.B0(In_Data[7]), 
	.A1(S_R_Data[7]), 
	.A0(n19));
   NOR3X2M U48 (.Y(n28), 
	.C(counter[1]), 
	.B(counter[3]), 
	.A(counter[2]));
   INVX2M U49 (.Y(n18), 
	.A(counter[0]));
   INVX2M U50 (.Y(n48), 
	.A(counter[1]));
endmodule

module FSM_test_1 (
	CLK, 
	RST, 
	Data_Valid, 
	PAR_EN, 
	ser_done, 
	mux_sel, 
	ser_en, 
	Basy, 
	Parity_Calc_En, 
	test_so, 
	test_se, 
	FE_OFN5_M_Domain2_SYNC_RST);
   input CLK;
   input RST;
   input Data_Valid;
   input PAR_EN;
   input ser_done;
   output [1:0] mux_sel;
   output ser_en;
   output Basy;
   output Parity_Calc_En;
   output test_so;
   input test_se;
   input FE_OFN5_M_Domain2_SYNC_RST;

   // Internal wires
   wire Basy_c;
   wire n8;
   wire n9;
   wire n10;
   wire n5;
   wire n6;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = current_state[2] ;
   assign Parity_Calc_En = next_state[1] ;

   SDFFRQX2M Basy_reg (.SI(ser_done), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Basy), 
	.D(Basy_c), 
	.CK(CLK));
   SDFFRQX2M \current_state_reg[0]  (.SI(Basy), 
	.SE(test_se), 
	.RN(RST), 
	.Q(current_state[0]), 
	.D(next_state[0]), 
	.CK(CLK));
   SDFFRQX2M \current_state_reg[1]  (.SI(n5), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(current_state[1]), 
	.D(next_state[1]), 
	.CK(CLK));
   SDFFRQX2M \current_state_reg[2]  (.SI(n6), 
	.SE(test_se), 
	.RN(RST), 
	.Q(current_state[2]), 
	.D(next_state[2]), 
	.CK(CLK));
   INVX2M U7 (.Y(mux_sel[0]), 
	.A(n10));
   NOR4X1M U8 (.Y(ser_en), 
	.D(n6), 
	.C(n5), 
	.B(current_state[2]), 
	.A(ser_done));
   NOR2X2M U9 (.Y(n10), 
	.B(current_state[2]), 
	.A(n5));
   AOI21X2M U10 (.Y(next_state[1]), 
	.B0(current_state[2]), 
	.A1(n5), 
	.A0(n6));
   OAI22X1M U11 (.Y(next_state[0]), 
	.B1(n9), 
	.B0(current_state[1]), 
	.A1(mux_sel[0]), 
	.A0(ser_done));
   AOI2B1X1M U12 (.Y(n9), 
	.B0(n10), 
	.A1N(current_state[2]), 
	.A0(Data_Valid));
   NOR2X2M U13 (.Y(mux_sel[1]), 
	.B(current_state[2]), 
	.A(n6));
   OAI21X2M U14 (.Y(Basy_c), 
	.B0(mux_sel[0]), 
	.A1(n6), 
	.A0(current_state[0]));
   INVX2M U15 (.Y(n5), 
	.A(current_state[0]));
   INVX2M U16 (.Y(n6), 
	.A(current_state[1]));
   NOR2BX2M U17 (.Y(next_state[2]), 
	.B(n8), 
	.AN(mux_sel[1]));
   AOI2B1X1M U18 (.Y(n8), 
	.B0(n5), 
	.A1N(PAR_EN), 
	.A0(ser_done));
endmodule

module UART_TOP_test_1 (
	CLK, 
	RST, 
	P_DATA, 
	Data_Valid, 
	PAR_EN, 
	PAR_TYP, 
	busy, 
	TX_OUT, 
	test_si2, 
	test_si1, 
	test_so1, 
	test_se, 
	FE_OFN5_M_Domain2_SYNC_RST, 
	TX_CLK_M__L3_N1, 
	TX_CLK_M__L3_N2, 
	TX_CLK_M__L3_N3);
   input CLK;
   input RST;
   input [7:0] P_DATA;
   input Data_Valid;
   input PAR_EN;
   input PAR_TYP;
   output busy;
   output TX_OUT;
   input test_si2;
   input test_si1;
   output test_so1;
   input test_se;
   input FE_OFN5_M_Domain2_SYNC_RST;
   input TX_CLK_M__L3_N1;
   input TX_CLK_M__L3_N2;
   input TX_CLK_M__L3_N3;

   // Internal wires
   wire ser_data;
   wire par_bit;
   wire Parity_Calc_En;
   wire ser_en;
   wire ser_done;
   wire [1:0] mux_sel;

   MUX_4x1_test_1 U1_MUX_4x1 (.CLK(CLK), 
	.RST(RST), 
	.mux_sel({ mux_sel[1],
		mux_sel[0] }), 
	.input_1(1'b0), 
	.input_2(1'b1), 
	.input_3(ser_data), 
	.input_4(par_bit), 
	.OUT(TX_OUT), 
	.test_si(test_si2), 
	.test_se(test_se));
   Parity_Calc_test_1 U2_Parity_Calc (.CLK(CLK), 
	.RST(RST), 
	.In_Data({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }), 
	.Data_Valid(Data_Valid), 
	.Basy_signal(busy), 
	.Parity_Calc_En(Parity_Calc_En), 
	.PAR_TYP(PAR_TYP), 
	.par_bit(par_bit), 
	.test_si(test_si1), 
	.test_se(test_se), 
	.TX_CLK_M__L3_N1(TX_CLK_M__L3_N1), 
	.TX_CLK_M__L3_N2(TX_CLK_M__L3_N2));
   Serializer_1byte_test_1 U3_Serializer (.In_Data({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }), 
	.Data_Valid(Data_Valid), 
	.Basy_signal(busy), 
	.CLK(CLK), 
	.RST(RST), 
	.ser_en(ser_en), 
	.ser_done(ser_done), 
	.Out_Data(ser_data), 
	.test_si(par_bit), 
	.test_se(test_se), 
	.FE_OFN5_M_Domain2_SYNC_RST(FE_OFN5_M_Domain2_SYNC_RST), 
	.TX_CLK_M__L3_N1(TX_CLK_M__L3_N1), 
	.TX_CLK_M__L3_N2(TX_CLK_M__L3_N2), 
	.TX_CLK_M__L3_N3(TX_CLK_M__L3_N3));
   FSM_test_1 U4_FSM (.CLK(CLK), 
	.RST(RST), 
	.Data_Valid(Data_Valid), 
	.PAR_EN(PAR_EN), 
	.ser_done(ser_done), 
	.mux_sel({ mux_sel[1],
		mux_sel[0] }), 
	.ser_en(ser_en), 
	.Basy(busy), 
	.Parity_Calc_En(Parity_Calc_En), 
	.test_so(test_so1), 
	.test_se(test_se), 
	.FE_OFN5_M_Domain2_SYNC_RST(FE_OFN5_M_Domain2_SYNC_RST));
endmodule

module FIFO_W_Addr_Size3_test_1 (
	W_CLK, 
	W_RST, 
	W_INC, 
	GR_Ptr_Syn, 
	FIFO_Full, 
	W_Addr, 
	GW_Ptr, 
	test_si, 
	test_se, 
	REF_CLK_M__L5_N5, 
	REF_CLK_M__L5_N6);
   input W_CLK;
   input W_RST;
   input W_INC;
   input [3:0] GR_Ptr_Syn;
   output FIFO_Full;
   output [2:0] W_Addr;
   output [3:0] GW_Ptr;
   input test_si;
   input test_se;
   input REF_CLK_M__L5_N5;
   input REF_CLK_M__L5_N6;

   // Internal wires
   wire \Address[3] ;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire [2:0] Comb_G_W_Ptr;

   SDFFRQX2M \Address_reg[3]  (.SI(W_Addr[2]), 
	.SE(test_se), 
	.RN(W_RST), 
	.Q(\Address[3] ), 
	.D(n19), 
	.CK(W_CLK));
   SDFFRQX2M \Address_reg[2]  (.SI(W_Addr[1]), 
	.SE(test_se), 
	.RN(W_RST), 
	.Q(W_Addr[2]), 
	.D(n20), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \GW_Ptr_reg[3]  (.SI(GW_Ptr[2]), 
	.SE(test_se), 
	.RN(W_RST), 
	.Q(GW_Ptr[3]), 
	.D(\Address[3] ), 
	.CK(W_CLK));
   SDFFRQX2M \GW_Ptr_reg[2]  (.SI(GW_Ptr[1]), 
	.SE(test_se), 
	.RN(W_RST), 
	.Q(GW_Ptr[2]), 
	.D(Comb_G_W_Ptr[2]), 
	.CK(W_CLK));
   SDFFRQX2M \GW_Ptr_reg[1]  (.SI(GW_Ptr[0]), 
	.SE(test_se), 
	.RN(W_RST), 
	.Q(GW_Ptr[1]), 
	.D(Comb_G_W_Ptr[1]), 
	.CK(W_CLK));
   SDFFRQX2M \GW_Ptr_reg[0]  (.SI(\Address[3] ), 
	.SE(test_se), 
	.RN(W_RST), 
	.Q(GW_Ptr[0]), 
	.D(Comb_G_W_Ptr[0]), 
	.CK(W_CLK));
   SDFFRQX2M \Address_reg[1]  (.SI(W_Addr[0]), 
	.SE(test_se), 
	.RN(W_RST), 
	.Q(W_Addr[1]), 
	.D(n21), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRX1M \Address_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(W_RST), 
	.QN(n9), 
	.Q(W_Addr[0]), 
	.D(n22), 
	.CK(REF_CLK_M__L5_N6));
   NAND2X2M U12 (.Y(n13), 
	.B(n14), 
	.A(W_INC));
   INVX2M U13 (.Y(FIFO_Full), 
	.A(n14));
   XNOR2X2M U14 (.Y(n15), 
	.B(GR_Ptr_Syn[1]), 
	.A(Comb_G_W_Ptr[1]));
   XNOR2X2M U15 (.Y(Comb_G_W_Ptr[0]), 
	.B(W_Addr[1]), 
	.A(n9));
   NOR2X2M U16 (.Y(n12), 
	.B(n9), 
	.A(n13));
   XNOR2X2M U17 (.Y(n20), 
	.B(n11), 
	.A(W_Addr[2]));
   XNOR2X2M U18 (.Y(n19), 
	.B(n10), 
	.A(\Address[3] ));
   NAND2BX2M U19 (.Y(n10), 
	.B(W_Addr[2]), 
	.AN(n11));
   NAND4X2M U20 (.Y(n14), 
	.D(n18), 
	.C(n17), 
	.B(n16), 
	.A(n15));
   CLKXOR2X2M U21 (.Y(n18), 
	.B(\Address[3] ), 
	.A(GR_Ptr_Syn[3]));
   XNOR2X2M U22 (.Y(n16), 
	.B(GR_Ptr_Syn[0]), 
	.A(Comb_G_W_Ptr[0]));
   CLKXOR2X2M U23 (.Y(n17), 
	.B(Comb_G_W_Ptr[2]), 
	.A(GR_Ptr_Syn[2]));
   NAND2X2M U24 (.Y(n11), 
	.B(W_Addr[1]), 
	.A(n12));
   CLKXOR2X2M U25 (.Y(Comb_G_W_Ptr[2]), 
	.B(W_Addr[2]), 
	.A(\Address[3] ));
   CLKXOR2X2M U26 (.Y(Comb_G_W_Ptr[1]), 
	.B(W_Addr[2]), 
	.A(W_Addr[1]));
   CLKXOR2X2M U27 (.Y(n21), 
	.B(n12), 
	.A(W_Addr[1]));
   CLKXOR2X2M U28 (.Y(n22), 
	.B(n13), 
	.A(n9));
endmodule

module BIT_SYNC_2_00000004_test_0 (
	CLK, 
	RST, 
	ASYNC, 
	SYNC, 
	test_se, 
	FE_OFN5_M_Domain2_SYNC_RST, 
	TX_CLK_M__L3_N3);
   input CLK;
   input RST;
   input [3:0] ASYNC;
   output [3:0] SYNC;
   input test_se;
   input FE_OFN5_M_Domain2_SYNC_RST;
   input TX_CLK_M__L3_N3;

   // Internal wires
   wire \sync_reg[3][0] ;
   wire \sync_reg[2][0] ;
   wire \sync_reg[1][0] ;
   wire \sync_reg[0][0] ;

   SDFFRQX2M \sync_reg_reg[2][1]  (.SI(\sync_reg[2][0] ), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(SYNC[2]), 
	.D(\sync_reg[2][0] ), 
	.CK(TX_CLK_M__L3_N3));
   SDFFRQX2M \sync_reg_reg[1][1]  (.SI(\sync_reg[1][0] ), 
	.SE(test_se), 
	.RN(RST), 
	.Q(SYNC[1]), 
	.D(\sync_reg[1][0] ), 
	.CK(CLK));
   SDFFRQX2M \sync_reg_reg[0][1]  (.SI(\sync_reg[0][0] ), 
	.SE(test_se), 
	.RN(RST), 
	.Q(SYNC[0]), 
	.D(\sync_reg[0][0] ), 
	.CK(CLK));
   SDFFRQX2M \sync_reg_reg[3][0]  (.SI(SYNC[2]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(\sync_reg[3][0] ), 
	.D(ASYNC[3]), 
	.CK(TX_CLK_M__L3_N3));
   SDFFRQX2M \sync_reg_reg[2][0]  (.SI(SYNC[1]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(\sync_reg[2][0] ), 
	.D(ASYNC[2]), 
	.CK(TX_CLK_M__L3_N3));
   SDFFRQX2M \sync_reg_reg[1][0]  (.SI(SYNC[0]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(\sync_reg[1][0] ), 
	.D(ASYNC[1]), 
	.CK(TX_CLK_M__L3_N3));
   SDFFRQX2M \sync_reg_reg[0][0]  (.SI(ASYNC[3]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(\sync_reg[0][0] ), 
	.D(ASYNC[0]), 
	.CK(CLK));
   SDFFRQX1M \sync_reg_reg[3][1]  (.SI(\sync_reg[3][0] ), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(SYNC[3]), 
	.D(\sync_reg[3][0] ), 
	.CK(TX_CLK_M__L3_N3));
endmodule

module FIFO_R_Addr_Size3_test_1 (
	R_CLK, 
	R_RST, 
	R_INC, 
	GW_Ptr_Syn, 
	FIFO_Empty, 
	R_Addr, 
	GR_Ptr, 
	test_se, 
	FE_OFN5_M_Domain2_SYNC_RST, 
	TX_CLK_M__L3_N3);
   input R_CLK;
   input R_RST;
   input R_INC;
   input [3:0] GW_Ptr_Syn;
   output FIFO_Empty;
   output [2:0] R_Addr;
   output [3:0] GR_Ptr;
   input test_se;
   input FE_OFN5_M_Domain2_SYNC_RST;
   input TX_CLK_M__L3_N3;

   // Internal wires
   wire \Address[3] ;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire [2:0] Comb_G_R_Ptr;

   SDFFRQX2M \Address_reg[3]  (.SI(R_Addr[2]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(\Address[3] ), 
	.D(n19), 
	.CK(TX_CLK_M__L3_N3));
   SDFFRX1M \Address_reg[0]  (.SI(GW_Ptr_Syn[3]), 
	.SE(test_se), 
	.RN(R_RST), 
	.QN(n9), 
	.Q(R_Addr[0]), 
	.D(n22), 
	.CK(TX_CLK_M__L3_N3));
   SDFFRQX2M \Address_reg[2]  (.SI(R_Addr[1]), 
	.SE(test_se), 
	.RN(R_RST), 
	.Q(R_Addr[2]), 
	.D(n20), 
	.CK(R_CLK));
   SDFFRQX2M \GR_Ptr_reg[3]  (.SI(GR_Ptr[2]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(GR_Ptr[3]), 
	.D(\Address[3] ), 
	.CK(TX_CLK_M__L3_N3));
   SDFFRQX2M \GR_Ptr_reg[2]  (.SI(GR_Ptr[1]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(GR_Ptr[2]), 
	.D(Comb_G_R_Ptr[2]), 
	.CK(TX_CLK_M__L3_N3));
   SDFFRQX2M \GR_Ptr_reg[1]  (.SI(GR_Ptr[0]), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(GR_Ptr[1]), 
	.D(Comb_G_R_Ptr[1]), 
	.CK(TX_CLK_M__L3_N3));
   SDFFRQX2M \GR_Ptr_reg[0]  (.SI(\Address[3] ), 
	.SE(test_se), 
	.RN(FE_OFN5_M_Domain2_SYNC_RST), 
	.Q(GR_Ptr[0]), 
	.D(Comb_G_R_Ptr[0]), 
	.CK(TX_CLK_M__L3_N3));
   SDFFRQX4M \Address_reg[1]  (.SI(R_Addr[0]), 
	.SE(test_se), 
	.RN(R_RST), 
	.Q(R_Addr[1]), 
	.D(n21), 
	.CK(R_CLK));
   XNOR2X2M U12 (.Y(n16), 
	.B(GW_Ptr_Syn[0]), 
	.A(Comb_G_R_Ptr[0]));
   XNOR2X2M U13 (.Y(Comb_G_R_Ptr[0]), 
	.B(R_Addr[1]), 
	.A(n9));
   NOR2X2M U14 (.Y(n12), 
	.B(n9), 
	.A(n13));
   XNOR2X2M U15 (.Y(n19), 
	.B(n10), 
	.A(\Address[3] ));
   NAND2BX2M U16 (.Y(n10), 
	.B(R_Addr[2]), 
	.AN(n11));
   NAND4X2M U17 (.Y(FIFO_Empty), 
	.D(n18), 
	.C(n17), 
	.B(n16), 
	.A(n15));
   XNOR2X2M U18 (.Y(n17), 
	.B(GW_Ptr_Syn[3]), 
	.A(\Address[3] ));
   XNOR2X2M U19 (.Y(n18), 
	.B(GW_Ptr_Syn[2]), 
	.A(Comb_G_R_Ptr[2]));
   XNOR2X2M U20 (.Y(n15), 
	.B(GW_Ptr_Syn[1]), 
	.A(Comb_G_R_Ptr[1]));
   NAND2X2M U21 (.Y(n11), 
	.B(R_Addr[1]), 
	.A(n12));
   NAND2X2M U22 (.Y(n13), 
	.B(FIFO_Empty), 
	.A(R_INC));
   CLKXOR2X2M U23 (.Y(Comb_G_R_Ptr[1]), 
	.B(R_Addr[2]), 
	.A(R_Addr[1]));
   CLKXOR2X2M U24 (.Y(Comb_G_R_Ptr[2]), 
	.B(R_Addr[2]), 
	.A(\Address[3] ));
   XNOR2X2M U25 (.Y(n20), 
	.B(n11), 
	.A(R_Addr[2]));
   CLKXOR2X2M U26 (.Y(n21), 
	.B(n12), 
	.A(R_Addr[1]));
   CLKXOR2X2M U27 (.Y(n22), 
	.B(n13), 
	.A(n9));
endmodule

module BIT_SYNC_2_00000004_test_1 (
	CLK, 
	RST, 
	ASYNC, 
	SYNC, 
	test_se);
   input CLK;
   input RST;
   input [3:0] ASYNC;
   output [3:0] SYNC;
   input test_se;

   // Internal wires
   wire \sync_reg[3][0] ;
   wire \sync_reg[2][0] ;
   wire \sync_reg[1][0] ;
   wire \sync_reg[0][0] ;

   SDFFRQX2M \sync_reg_reg[1][1]  (.SI(\sync_reg[1][0] ), 
	.SE(test_se), 
	.RN(RST), 
	.Q(SYNC[1]), 
	.D(\sync_reg[1][0] ), 
	.CK(CLK));
   SDFFRQX2M \sync_reg_reg[0][1]  (.SI(\sync_reg[0][0] ), 
	.SE(test_se), 
	.RN(RST), 
	.Q(SYNC[0]), 
	.D(\sync_reg[0][0] ), 
	.CK(CLK));
   SDFFRQX2M \sync_reg_reg[3][1]  (.SI(\sync_reg[3][0] ), 
	.SE(test_se), 
	.RN(RST), 
	.Q(SYNC[3]), 
	.D(\sync_reg[3][0] ), 
	.CK(CLK));
   SDFFRQX2M \sync_reg_reg[2][1]  (.SI(\sync_reg[2][0] ), 
	.SE(test_se), 
	.RN(RST), 
	.Q(SYNC[2]), 
	.D(\sync_reg[2][0] ), 
	.CK(CLK));
   SDFFRQX2M \sync_reg_reg[3][0]  (.SI(SYNC[2]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(\sync_reg[3][0] ), 
	.D(ASYNC[3]), 
	.CK(CLK));
   SDFFRQX2M \sync_reg_reg[2][0]  (.SI(SYNC[1]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(\sync_reg[2][0] ), 
	.D(ASYNC[2]), 
	.CK(CLK));
   SDFFRQX2M \sync_reg_reg[1][0]  (.SI(SYNC[0]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(\sync_reg[1][0] ), 
	.D(ASYNC[1]), 
	.CK(CLK));
   SDFFRQX2M \sync_reg_reg[0][0]  (.SI(ASYNC[3]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(\sync_reg[0][0] ), 
	.D(ASYNC[0]), 
	.CK(CLK));
endmodule

module FIFO_MEM_Data_Width8_Addr_Size3_FIFO_Dipth8_test_1 (
	W_CLK, 
	W_RST, 
	W_INC, 
	FIFO_Full, 
	W_Addr, 
	W_Data, 
	R_Addr, 
	R_Data, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN1_M_Domain1_SYNC_RST, 
	FE_OFN4_M_Domain1_SYNC_RST, 
	REF_CLK_M__L5_N1, 
	REF_CLK_M__L5_N4, 
	REF_CLK_M__L5_N5, 
	REF_CLK_M__L5_N6, 
	REF_CLK_M__L5_N7);
   input W_CLK;
   input W_RST;
   input W_INC;
   input FIFO_Full;
   input [2:0] W_Addr;
   input [7:0] W_Data;
   input [2:0] R_Addr;
   output [7:0] R_Data;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN1_M_Domain1_SYNC_RST;
   input FE_OFN4_M_Domain1_SYNC_RST;
   input REF_CLK_M__L5_N1;
   input REF_CLK_M__L5_N4;
   input REF_CLK_M__L5_N5;
   input REF_CLK_M__L5_N6;
   input REF_CLK_M__L5_N7;

   // Internal wires
   wire N9;
   wire N10;
   wire N11;
   wire \memory[0][7] ;
   wire \memory[0][6] ;
   wire \memory[0][5] ;
   wire \memory[0][4] ;
   wire \memory[0][3] ;
   wire \memory[0][2] ;
   wire \memory[0][1] ;
   wire \memory[0][0] ;
   wire \memory[1][7] ;
   wire \memory[1][6] ;
   wire \memory[1][5] ;
   wire \memory[1][4] ;
   wire \memory[1][3] ;
   wire \memory[1][2] ;
   wire \memory[1][1] ;
   wire \memory[1][0] ;
   wire \memory[2][7] ;
   wire \memory[2][6] ;
   wire \memory[2][5] ;
   wire \memory[2][4] ;
   wire \memory[2][3] ;
   wire \memory[2][2] ;
   wire \memory[2][1] ;
   wire \memory[2][0] ;
   wire \memory[3][7] ;
   wire \memory[3][6] ;
   wire \memory[3][5] ;
   wire \memory[3][4] ;
   wire \memory[3][3] ;
   wire \memory[3][2] ;
   wire \memory[3][1] ;
   wire \memory[3][0] ;
   wire \memory[4][7] ;
   wire \memory[4][6] ;
   wire \memory[4][5] ;
   wire \memory[4][4] ;
   wire \memory[4][3] ;
   wire \memory[4][2] ;
   wire \memory[4][1] ;
   wire \memory[4][0] ;
   wire \memory[5][7] ;
   wire \memory[5][6] ;
   wire \memory[5][5] ;
   wire \memory[5][4] ;
   wire \memory[5][3] ;
   wire \memory[5][2] ;
   wire \memory[5][1] ;
   wire \memory[5][0] ;
   wire \memory[6][7] ;
   wire \memory[6][6] ;
   wire \memory[6][5] ;
   wire \memory[6][4] ;
   wire \memory[6][3] ;
   wire \memory[6][2] ;
   wire \memory[6][1] ;
   wire \memory[6][0] ;
   wire \memory[7][7] ;
   wire \memory[7][6] ;
   wire \memory[7][5] ;
   wire \memory[7][4] ;
   wire \memory[7][3] ;
   wire \memory[7][2] ;
   wire \memory[7][1] ;
   wire \memory[7][0] ;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;

   assign N9 = R_Addr[0] ;
   assign N10 = R_Addr[1] ;
   assign N11 = R_Addr[2] ;
   assign test_so1 = \memory[6][1]  ;
   assign test_so2 = \memory[7][7]  ;

   SDFFRQX2M \memory_reg[1][7]  (.SI(\memory[1][6] ), 
	.SE(n188), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[1][7] ), 
	.D(n141), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \memory_reg[1][6]  (.SI(\memory[1][5] ), 
	.SE(n187), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[1][6] ), 
	.D(n140), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[1][5]  (.SI(\memory[1][4] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[1][5] ), 
	.D(n139), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[1][4]  (.SI(\memory[1][3] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[1][4] ), 
	.D(n138), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[1][3]  (.SI(\memory[1][2] ), 
	.SE(n188), 
	.RN(W_RST), 
	.Q(\memory[1][3] ), 
	.D(n137), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[1][2]  (.SI(\memory[1][1] ), 
	.SE(n187), 
	.RN(W_RST), 
	.Q(\memory[1][2] ), 
	.D(n136), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[1][1]  (.SI(\memory[1][0] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[1][1] ), 
	.D(n135), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[1][0]  (.SI(\memory[0][7] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[1][0] ), 
	.D(n134), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[5][7]  (.SI(\memory[5][6] ), 
	.SE(n188), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[5][7] ), 
	.D(n109), 
	.CK(W_CLK));
   SDFFRQX2M \memory_reg[5][6]  (.SI(\memory[5][5] ), 
	.SE(n187), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[5][6] ), 
	.D(n108), 
	.CK(W_CLK));
   SDFFRQX2M \memory_reg[5][5]  (.SI(\memory[5][4] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[5][5] ), 
	.D(n107), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[5][4]  (.SI(\memory[5][3] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[5][4] ), 
	.D(n106), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[5][3]  (.SI(\memory[5][2] ), 
	.SE(n188), 
	.RN(W_RST), 
	.Q(\memory[5][3] ), 
	.D(n105), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[5][2]  (.SI(\memory[5][1] ), 
	.SE(n187), 
	.RN(W_RST), 
	.Q(\memory[5][2] ), 
	.D(n104), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[5][1]  (.SI(\memory[5][0] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[5][1] ), 
	.D(n103), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[5][0]  (.SI(\memory[4][7] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[5][0] ), 
	.D(n102), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[3][7]  (.SI(\memory[3][6] ), 
	.SE(n188), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[3][7] ), 
	.D(n125), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \memory_reg[3][6]  (.SI(\memory[3][5] ), 
	.SE(n187), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(\memory[3][6] ), 
	.D(n124), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \memory_reg[3][5]  (.SI(\memory[3][4] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[3][5] ), 
	.D(n123), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[3][4]  (.SI(\memory[3][3] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[3][4] ), 
	.D(n122), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[3][3]  (.SI(\memory[3][2] ), 
	.SE(n188), 
	.RN(W_RST), 
	.Q(\memory[3][3] ), 
	.D(n121), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[3][2]  (.SI(\memory[3][1] ), 
	.SE(n187), 
	.RN(W_RST), 
	.Q(\memory[3][2] ), 
	.D(n120), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[3][1]  (.SI(\memory[3][0] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[3][1] ), 
	.D(n119), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[3][0]  (.SI(\memory[2][7] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[3][0] ), 
	.D(n118), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[7][7]  (.SI(\memory[7][6] ), 
	.SE(n188), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[7][7] ), 
	.D(n93), 
	.CK(W_CLK));
   SDFFRQX2M \memory_reg[7][6]  (.SI(\memory[7][5] ), 
	.SE(n187), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[7][6] ), 
	.D(n92), 
	.CK(W_CLK));
   SDFFRQX2M \memory_reg[7][5]  (.SI(\memory[7][4] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[7][5] ), 
	.D(n91), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[7][4]  (.SI(\memory[7][3] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[7][4] ), 
	.D(n90), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[7][3]  (.SI(\memory[7][2] ), 
	.SE(n188), 
	.RN(W_RST), 
	.Q(\memory[7][3] ), 
	.D(n89), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \memory_reg[7][2]  (.SI(\memory[7][1] ), 
	.SE(n187), 
	.RN(W_RST), 
	.Q(\memory[7][2] ), 
	.D(n88), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[7][1]  (.SI(\memory[7][0] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[7][1] ), 
	.D(n87), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[7][0]  (.SI(\memory[6][7] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[7][0] ), 
	.D(n86), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[2][7]  (.SI(\memory[2][6] ), 
	.SE(n188), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[2][7] ), 
	.D(n133), 
	.CK(W_CLK));
   SDFFRQX2M \memory_reg[2][6]  (.SI(\memory[2][5] ), 
	.SE(n187), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[2][6] ), 
	.D(n132), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \memory_reg[2][5]  (.SI(\memory[2][4] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[2][5] ), 
	.D(n131), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[2][4]  (.SI(\memory[2][3] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[2][4] ), 
	.D(n130), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[2][3]  (.SI(\memory[2][2] ), 
	.SE(n188), 
	.RN(W_RST), 
	.Q(\memory[2][3] ), 
	.D(n129), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[2][2]  (.SI(\memory[2][1] ), 
	.SE(n187), 
	.RN(W_RST), 
	.Q(\memory[2][2] ), 
	.D(n128), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[2][1]  (.SI(\memory[2][0] ), 
	.SE(n186), 
	.RN(W_RST), 
	.Q(\memory[2][1] ), 
	.D(n127), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[2][0]  (.SI(\memory[1][7] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[2][0] ), 
	.D(n126), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[6][7]  (.SI(\memory[6][6] ), 
	.SE(n188), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[6][7] ), 
	.D(n101), 
	.CK(W_CLK));
   SDFFRQX2M \memory_reg[6][6]  (.SI(\memory[6][5] ), 
	.SE(n187), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[6][6] ), 
	.D(n100), 
	.CK(W_CLK));
   SDFFRQX2M \memory_reg[6][5]  (.SI(\memory[6][4] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[6][5] ), 
	.D(n99), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[6][4]  (.SI(\memory[6][3] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[6][4] ), 
	.D(n98), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \memory_reg[6][3]  (.SI(\memory[6][2] ), 
	.SE(n188), 
	.RN(W_RST), 
	.Q(\memory[6][3] ), 
	.D(n97), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \memory_reg[6][2]  (.SI(test_si2), 
	.SE(n187), 
	.RN(W_RST), 
	.Q(\memory[6][2] ), 
	.D(n96), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX4M \memory_reg[6][1]  (.SI(\memory[6][0] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[6][1] ), 
	.D(n95), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[6][0]  (.SI(\memory[5][7] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[6][0] ), 
	.D(n94), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[0][7]  (.SI(\memory[0][6] ), 
	.SE(n188), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[0][7] ), 
	.D(n149), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \memory_reg[0][6]  (.SI(\memory[0][5] ), 
	.SE(n187), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[0][6] ), 
	.D(n148), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \memory_reg[0][5]  (.SI(\memory[0][4] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[0][5] ), 
	.D(n147), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[0][4]  (.SI(\memory[0][3] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[0][4] ), 
	.D(n146), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[0][3]  (.SI(\memory[0][2] ), 
	.SE(n188), 
	.RN(W_RST), 
	.Q(\memory[0][3] ), 
	.D(n145), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[0][2]  (.SI(\memory[0][1] ), 
	.SE(n187), 
	.RN(W_RST), 
	.Q(\memory[0][2] ), 
	.D(n144), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[0][1]  (.SI(\memory[0][0] ), 
	.SE(n186), 
	.RN(W_RST), 
	.Q(\memory[0][1] ), 
	.D(n143), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[0][0]  (.SI(test_si1), 
	.SE(n185), 
	.RN(W_RST), 
	.Q(\memory[0][0] ), 
	.D(n142), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[4][7]  (.SI(\memory[4][6] ), 
	.SE(n188), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[4][7] ), 
	.D(n117), 
	.CK(W_CLK));
   SDFFRQX2M \memory_reg[4][6]  (.SI(\memory[4][5] ), 
	.SE(n187), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[4][6] ), 
	.D(n116), 
	.CK(W_CLK));
   SDFFRQX2M \memory_reg[4][5]  (.SI(\memory[4][4] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[4][5] ), 
	.D(n115), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[4][4]  (.SI(\memory[4][3] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[4][4] ), 
	.D(n114), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[4][3]  (.SI(\memory[4][2] ), 
	.SE(n188), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[4][3] ), 
	.D(n113), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \memory_reg[4][2]  (.SI(\memory[4][1] ), 
	.SE(n187), 
	.RN(W_RST), 
	.Q(\memory[4][2] ), 
	.D(n112), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \memory_reg[4][1]  (.SI(\memory[4][0] ), 
	.SE(n186), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[4][1] ), 
	.D(n111), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \memory_reg[4][0]  (.SI(\memory[3][7] ), 
	.SE(n185), 
	.RN(FE_OFN1_M_Domain1_SYNC_RST), 
	.Q(\memory[4][0] ), 
	.D(n110), 
	.CK(REF_CLK_M__L5_N7));
   NOR2BX2M U78 (.Y(n80), 
	.B(FIFO_Full), 
	.AN(W_INC));
   NAND3X2M U81 (.Y(n79), 
	.C(n76), 
	.B(n180), 
	.A(n179));
   NAND3X2M U82 (.Y(n85), 
	.C(n82), 
	.B(n180), 
	.A(n179));
   NOR2BX2M U83 (.Y(n82), 
	.B(W_Addr[2]), 
	.AN(n80));
   OAI2BB2X1M U84 (.Y(n142), 
	.B1(n85), 
	.B0(n178), 
	.A1N(n85), 
	.A0N(\memory[0][0] ));
   OAI2BB2X1M U85 (.Y(n143), 
	.B1(n85), 
	.B0(n177), 
	.A1N(n85), 
	.A0N(\memory[0][1] ));
   OAI2BB2X1M U86 (.Y(n144), 
	.B1(n85), 
	.B0(n176), 
	.A1N(n85), 
	.A0N(\memory[0][2] ));
   OAI2BB2X1M U87 (.Y(n145), 
	.B1(n85), 
	.B0(n175), 
	.A1N(n85), 
	.A0N(\memory[0][3] ));
   OAI2BB2X1M U88 (.Y(n146), 
	.B1(n85), 
	.B0(n174), 
	.A1N(n85), 
	.A0N(\memory[0][4] ));
   OAI2BB2X1M U89 (.Y(n147), 
	.B1(n85), 
	.B0(n173), 
	.A1N(n85), 
	.A0N(\memory[0][5] ));
   OAI2BB2X1M U90 (.Y(n148), 
	.B1(n85), 
	.B0(n172), 
	.A1N(n85), 
	.A0N(\memory[0][6] ));
   OAI2BB2X1M U91 (.Y(n149), 
	.B1(n85), 
	.B0(n171), 
	.A1N(n85), 
	.A0N(\memory[0][7] ));
   OAI2BB2X1M U92 (.Y(n110), 
	.B1(n79), 
	.B0(n178), 
	.A1N(n79), 
	.A0N(\memory[4][0] ));
   OAI2BB2X1M U93 (.Y(n111), 
	.B1(n79), 
	.B0(n177), 
	.A1N(n79), 
	.A0N(\memory[4][1] ));
   OAI2BB2X1M U94 (.Y(n112), 
	.B1(n79), 
	.B0(n176), 
	.A1N(n79), 
	.A0N(\memory[4][2] ));
   OAI2BB2X1M U95 (.Y(n113), 
	.B1(n79), 
	.B0(n175), 
	.A1N(n79), 
	.A0N(\memory[4][3] ));
   OAI2BB2X1M U96 (.Y(n114), 
	.B1(n79), 
	.B0(n174), 
	.A1N(n79), 
	.A0N(\memory[4][4] ));
   OAI2BB2X1M U97 (.Y(n115), 
	.B1(n79), 
	.B0(n173), 
	.A1N(n79), 
	.A0N(\memory[4][5] ));
   OAI2BB2X1M U98 (.Y(n116), 
	.B1(n79), 
	.B0(n172), 
	.A1N(n79), 
	.A0N(\memory[4][6] ));
   OAI2BB2X1M U99 (.Y(n117), 
	.B1(n79), 
	.B0(n171), 
	.A1N(n79), 
	.A0N(\memory[4][7] ));
   INVX2M U100 (.Y(n178), 
	.A(W_Data[0]));
   INVX2M U101 (.Y(n177), 
	.A(W_Data[1]));
   INVX2M U102 (.Y(n176), 
	.A(W_Data[2]));
   INVX2M U103 (.Y(n175), 
	.A(W_Data[3]));
   INVX2M U104 (.Y(n174), 
	.A(W_Data[4]));
   INVX2M U105 (.Y(n173), 
	.A(W_Data[5]));
   INVX2M U106 (.Y(n172), 
	.A(W_Data[6]));
   INVX2M U107 (.Y(n171), 
	.A(W_Data[7]));
   OAI2BB2X1M U108 (.Y(n94), 
	.B1(n77), 
	.B0(n178), 
	.A1N(n77), 
	.A0N(\memory[6][0] ));
   OAI2BB2X1M U109 (.Y(n95), 
	.B1(n77), 
	.B0(n177), 
	.A1N(n77), 
	.A0N(\memory[6][1] ));
   OAI2BB2X1M U110 (.Y(n96), 
	.B1(n77), 
	.B0(n176), 
	.A1N(n77), 
	.A0N(\memory[6][2] ));
   OAI2BB2X1M U111 (.Y(n97), 
	.B1(n77), 
	.B0(n175), 
	.A1N(n77), 
	.A0N(\memory[6][3] ));
   OAI2BB2X1M U112 (.Y(n98), 
	.B1(n77), 
	.B0(n174), 
	.A1N(n77), 
	.A0N(\memory[6][4] ));
   OAI2BB2X1M U113 (.Y(n99), 
	.B1(n77), 
	.B0(n173), 
	.A1N(n77), 
	.A0N(\memory[6][5] ));
   OAI2BB2X1M U114 (.Y(n100), 
	.B1(n77), 
	.B0(n172), 
	.A1N(n77), 
	.A0N(\memory[6][6] ));
   OAI2BB2X1M U115 (.Y(n101), 
	.B1(n77), 
	.B0(n171), 
	.A1N(n77), 
	.A0N(\memory[6][7] ));
   OAI2BB2X1M U116 (.Y(n102), 
	.B1(n78), 
	.B0(n178), 
	.A1N(n78), 
	.A0N(\memory[5][0] ));
   OAI2BB2X1M U117 (.Y(n103), 
	.B1(n78), 
	.B0(n177), 
	.A1N(n78), 
	.A0N(\memory[5][1] ));
   OAI2BB2X1M U118 (.Y(n104), 
	.B1(n78), 
	.B0(n176), 
	.A1N(n78), 
	.A0N(\memory[5][2] ));
   OAI2BB2X1M U119 (.Y(n105), 
	.B1(n78), 
	.B0(n175), 
	.A1N(n78), 
	.A0N(\memory[5][3] ));
   OAI2BB2X1M U120 (.Y(n106), 
	.B1(n78), 
	.B0(n174), 
	.A1N(n78), 
	.A0N(\memory[5][4] ));
   OAI2BB2X1M U121 (.Y(n107), 
	.B1(n78), 
	.B0(n173), 
	.A1N(n78), 
	.A0N(\memory[5][5] ));
   OAI2BB2X1M U122 (.Y(n108), 
	.B1(n78), 
	.B0(n172), 
	.A1N(n78), 
	.A0N(\memory[5][6] ));
   OAI2BB2X1M U123 (.Y(n109), 
	.B1(n78), 
	.B0(n171), 
	.A1N(n78), 
	.A0N(\memory[5][7] ));
   OAI2BB2X1M U124 (.Y(n118), 
	.B1(n81), 
	.B0(n178), 
	.A1N(n81), 
	.A0N(\memory[3][0] ));
   OAI2BB2X1M U125 (.Y(n119), 
	.B1(n81), 
	.B0(n177), 
	.A1N(n81), 
	.A0N(\memory[3][1] ));
   OAI2BB2X1M U126 (.Y(n120), 
	.B1(n81), 
	.B0(n176), 
	.A1N(n81), 
	.A0N(\memory[3][2] ));
   OAI2BB2X1M U127 (.Y(n121), 
	.B1(n81), 
	.B0(n175), 
	.A1N(n81), 
	.A0N(\memory[3][3] ));
   OAI2BB2X1M U128 (.Y(n122), 
	.B1(n81), 
	.B0(n174), 
	.A1N(n81), 
	.A0N(\memory[3][4] ));
   OAI2BB2X1M U129 (.Y(n123), 
	.B1(n81), 
	.B0(n173), 
	.A1N(n81), 
	.A0N(\memory[3][5] ));
   OAI2BB2X1M U130 (.Y(n124), 
	.B1(n81), 
	.B0(n172), 
	.A1N(n81), 
	.A0N(\memory[3][6] ));
   OAI2BB2X1M U131 (.Y(n125), 
	.B1(n81), 
	.B0(n171), 
	.A1N(n81), 
	.A0N(\memory[3][7] ));
   OAI2BB2X1M U132 (.Y(n126), 
	.B1(n83), 
	.B0(n178), 
	.A1N(n83), 
	.A0N(\memory[2][0] ));
   OAI2BB2X1M U133 (.Y(n127), 
	.B1(n83), 
	.B0(n177), 
	.A1N(n83), 
	.A0N(\memory[2][1] ));
   OAI2BB2X1M U134 (.Y(n128), 
	.B1(n83), 
	.B0(n176), 
	.A1N(n83), 
	.A0N(\memory[2][2] ));
   OAI2BB2X1M U135 (.Y(n129), 
	.B1(n83), 
	.B0(n175), 
	.A1N(n83), 
	.A0N(\memory[2][3] ));
   OAI2BB2X1M U136 (.Y(n130), 
	.B1(n83), 
	.B0(n174), 
	.A1N(n83), 
	.A0N(\memory[2][4] ));
   OAI2BB2X1M U137 (.Y(n131), 
	.B1(n83), 
	.B0(n173), 
	.A1N(n83), 
	.A0N(\memory[2][5] ));
   OAI2BB2X1M U138 (.Y(n132), 
	.B1(n83), 
	.B0(n172), 
	.A1N(n83), 
	.A0N(\memory[2][6] ));
   OAI2BB2X1M U139 (.Y(n133), 
	.B1(n83), 
	.B0(n171), 
	.A1N(n83), 
	.A0N(\memory[2][7] ));
   OAI2BB2X1M U140 (.Y(n134), 
	.B1(n84), 
	.B0(n178), 
	.A1N(n84), 
	.A0N(\memory[1][0] ));
   OAI2BB2X1M U141 (.Y(n135), 
	.B1(n84), 
	.B0(n177), 
	.A1N(n84), 
	.A0N(\memory[1][1] ));
   OAI2BB2X1M U142 (.Y(n136), 
	.B1(n84), 
	.B0(n176), 
	.A1N(n84), 
	.A0N(\memory[1][2] ));
   OAI2BB2X1M U143 (.Y(n137), 
	.B1(n84), 
	.B0(n175), 
	.A1N(n84), 
	.A0N(\memory[1][3] ));
   OAI2BB2X1M U144 (.Y(n138), 
	.B1(n84), 
	.B0(n174), 
	.A1N(n84), 
	.A0N(\memory[1][4] ));
   OAI2BB2X1M U145 (.Y(n139), 
	.B1(n84), 
	.B0(n173), 
	.A1N(n84), 
	.A0N(\memory[1][5] ));
   OAI2BB2X1M U146 (.Y(n140), 
	.B1(n84), 
	.B0(n172), 
	.A1N(n84), 
	.A0N(\memory[1][6] ));
   OAI2BB2X1M U147 (.Y(n141), 
	.B1(n84), 
	.B0(n171), 
	.A1N(n84), 
	.A0N(\memory[1][7] ));
   OAI2BB2X1M U148 (.Y(n86), 
	.B1(n178), 
	.B0(n75), 
	.A1N(n75), 
	.A0N(\memory[7][0] ));
   OAI2BB2X1M U149 (.Y(n87), 
	.B1(n177), 
	.B0(n75), 
	.A1N(n75), 
	.A0N(\memory[7][1] ));
   OAI2BB2X1M U150 (.Y(n88), 
	.B1(n176), 
	.B0(n75), 
	.A1N(n75), 
	.A0N(\memory[7][2] ));
   OAI2BB2X1M U151 (.Y(n89), 
	.B1(n175), 
	.B0(n75), 
	.A1N(n75), 
	.A0N(\memory[7][3] ));
   OAI2BB2X1M U152 (.Y(n90), 
	.B1(n174), 
	.B0(n75), 
	.A1N(n75), 
	.A0N(\memory[7][4] ));
   OAI2BB2X1M U153 (.Y(n91), 
	.B1(n173), 
	.B0(n75), 
	.A1N(n75), 
	.A0N(\memory[7][5] ));
   OAI2BB2X1M U154 (.Y(n92), 
	.B1(n172), 
	.B0(n75), 
	.A1N(n75), 
	.A0N(\memory[7][6] ));
   OAI2BB2X1M U155 (.Y(n93), 
	.B1(n171), 
	.B0(n75), 
	.A1N(n75), 
	.A0N(\memory[7][7] ));
   AND2X2M U156 (.Y(n76), 
	.B(n80), 
	.A(W_Addr[2]));
   NAND3X2M U157 (.Y(n78), 
	.C(W_Addr[0]), 
	.B(n180), 
	.A(n76));
   NAND3X2M U158 (.Y(n81), 
	.C(n82), 
	.B(W_Addr[0]), 
	.A(W_Addr[1]));
   NAND3X2M U159 (.Y(n84), 
	.C(n82), 
	.B(n180), 
	.A(W_Addr[0]));
   NAND3X2M U160 (.Y(n83), 
	.C(n82), 
	.B(n179), 
	.A(W_Addr[1]));
   NAND3X2M U161 (.Y(n75), 
	.C(W_Addr[1]), 
	.B(n76), 
	.A(W_Addr[0]));
   NAND3X2M U162 (.Y(n77), 
	.C(W_Addr[1]), 
	.B(n179), 
	.A(n76));
   INVX2M U163 (.Y(n179), 
	.A(W_Addr[0]));
   INVX2M U164 (.Y(n180), 
	.A(W_Addr[1]));
   BUFX4M U165 (.Y(n156), 
	.A(N9));
   MX2X2M U166 (.Y(R_Data[7]), 
	.S0(N11), 
	.B(n154), 
	.A(n155));
   MX4X1M U167 (.Y(n155), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[3][7] ), 
	.C(\memory[2][7] ), 
	.B(\memory[1][7] ), 
	.A(\memory[0][7] ));
   MX4X1M U168 (.Y(n154), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[7][7] ), 
	.C(\memory[6][7] ), 
	.B(\memory[5][7] ), 
	.A(\memory[4][7] ));
   MX2X2M U169 (.Y(R_Data[0]), 
	.S0(N11), 
	.B(n65), 
	.A(n66));
   MX4X1M U170 (.Y(n66), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[3][0] ), 
	.C(\memory[2][0] ), 
	.B(\memory[1][0] ), 
	.A(\memory[0][0] ));
   MX4X1M U171 (.Y(n65), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[7][0] ), 
	.C(\memory[6][0] ), 
	.B(\memory[5][0] ), 
	.A(\memory[4][0] ));
   MX2X2M U172 (.Y(R_Data[1]), 
	.S0(N11), 
	.B(n67), 
	.A(n68));
   MX4X1M U173 (.Y(n68), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[3][1] ), 
	.C(\memory[2][1] ), 
	.B(\memory[1][1] ), 
	.A(\memory[0][1] ));
   MX4X1M U174 (.Y(n67), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[7][1] ), 
	.C(\memory[6][1] ), 
	.B(\memory[5][1] ), 
	.A(\memory[4][1] ));
   MX2X2M U175 (.Y(R_Data[2]), 
	.S0(N11), 
	.B(n69), 
	.A(n70));
   MX4X1M U176 (.Y(n70), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[3][2] ), 
	.C(\memory[2][2] ), 
	.B(\memory[1][2] ), 
	.A(\memory[0][2] ));
   MX4X1M U177 (.Y(n69), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[7][2] ), 
	.C(\memory[6][2] ), 
	.B(\memory[5][2] ), 
	.A(\memory[4][2] ));
   MX2X2M U178 (.Y(R_Data[3]), 
	.S0(N11), 
	.B(n71), 
	.A(n72));
   MX4X1M U179 (.Y(n72), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[3][3] ), 
	.C(\memory[2][3] ), 
	.B(\memory[1][3] ), 
	.A(\memory[0][3] ));
   MX4X1M U180 (.Y(n71), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[7][3] ), 
	.C(\memory[6][3] ), 
	.B(\memory[5][3] ), 
	.A(\memory[4][3] ));
   MX2X2M U181 (.Y(R_Data[4]), 
	.S0(N11), 
	.B(n73), 
	.A(n74));
   MX4X1M U182 (.Y(n74), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[3][4] ), 
	.C(\memory[2][4] ), 
	.B(\memory[1][4] ), 
	.A(\memory[0][4] ));
   MX4X1M U183 (.Y(n73), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[7][4] ), 
	.C(\memory[6][4] ), 
	.B(\memory[5][4] ), 
	.A(\memory[4][4] ));
   MX2X2M U184 (.Y(R_Data[5]), 
	.S0(N11), 
	.B(n150), 
	.A(n151));
   MX4X1M U185 (.Y(n151), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[3][5] ), 
	.C(\memory[2][5] ), 
	.B(\memory[1][5] ), 
	.A(\memory[0][5] ));
   MX4X1M U186 (.Y(n150), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[7][5] ), 
	.C(\memory[6][5] ), 
	.B(\memory[5][5] ), 
	.A(\memory[4][5] ));
   MX2X2M U187 (.Y(R_Data[6]), 
	.S0(N11), 
	.B(n152), 
	.A(n153));
   MX4X1M U188 (.Y(n153), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[3][6] ), 
	.C(\memory[2][6] ), 
	.B(\memory[1][6] ), 
	.A(\memory[0][6] ));
   MX4X1M U189 (.Y(n152), 
	.S1(N10), 
	.S0(n156), 
	.D(\memory[7][6] ), 
	.C(\memory[6][6] ), 
	.B(\memory[5][6] ), 
	.A(\memory[4][6] ));
   INVXLM U190 (.Y(n184), 
	.A(test_se));
   CLKINVX2M U191 (.Y(n185), 
	.A(n184));
   CLKINVX2M U192 (.Y(n186), 
	.A(n184));
   CLKINVX2M U193 (.Y(n187), 
	.A(n184));
   CLKINVX2M U194 (.Y(n188), 
	.A(n184));
endmodule

module AS_FIFO_TOP_Data_Width8_Addr_Size3_FIFO_Dipth8_NUM_STAGES2_test_1 (
	I_W_CLK, 
	I_W_RST, 
	I_W_INC, 
	I_Data, 
	I_R_CLK, 
	I_R_RST, 
	I_R_INC, 
	O_Data, 
	FIFO_Full, 
	FIFO_Empty, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN1_M_Domain1_SYNC_RST, 
	FE_OFN4_M_Domain1_SYNC_RST, 
	FE_OFN5_M_Domain2_SYNC_RST, 
	TX_CLK_M__L3_N3, 
	REF_CLK_M__L5_N1, 
	REF_CLK_M__L5_N4, 
	REF_CLK_M__L5_N5, 
	REF_CLK_M__L5_N6, 
	REF_CLK_M__L5_N7);
   input I_W_CLK;
   input I_W_RST;
   input I_W_INC;
   input [7:0] I_Data;
   input I_R_CLK;
   input I_R_RST;
   input I_R_INC;
   output [7:0] O_Data;
   output FIFO_Full;
   output FIFO_Empty;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN1_M_Domain1_SYNC_RST;
   input FE_OFN4_M_Domain1_SYNC_RST;
   input FE_OFN5_M_Domain2_SYNC_RST;
   input TX_CLK_M__L3_N3;
   input REF_CLK_M__L5_N1;
   input REF_CLK_M__L5_N4;
   input REF_CLK_M__L5_N5;
   input REF_CLK_M__L5_N6;
   input REF_CLK_M__L5_N7;

   // Internal wires
   wire [3:0] GR_Ptr_Syn;
   wire [2:0] W_Addr;
   wire [3:0] GW_Ptr;
   wire [3:0] GW_Ptr_Syn;
   wire [2:0] R_Addr;
   wire [3:0] GR_Ptr;

   FIFO_W_Addr_Size3_test_1 U0_FIFO_W (.W_CLK(REF_CLK_M__L5_N4), 
	.W_RST(I_W_RST), 
	.W_INC(I_W_INC), 
	.GR_Ptr_Syn({ GR_Ptr_Syn[3],
		GR_Ptr_Syn[2],
		GR_Ptr_Syn[1],
		GR_Ptr_Syn[0] }), 
	.FIFO_Full(FIFO_Full), 
	.W_Addr({ W_Addr[2],
		W_Addr[1],
		W_Addr[0] }), 
	.GW_Ptr({ GW_Ptr[3],
		GW_Ptr[2],
		GW_Ptr[1],
		GW_Ptr[0] }), 
	.test_si(test_si1), 
	.test_se(test_se), 
	.REF_CLK_M__L5_N5(REF_CLK_M__L5_N5), 
	.REF_CLK_M__L5_N6(REF_CLK_M__L5_N6));
   BIT_SYNC_2_00000004_test_0 U1_W2R_SYNC (.CLK(I_R_CLK), 
	.RST(I_R_RST), 
	.ASYNC({ GW_Ptr[3],
		GW_Ptr[2],
		GW_Ptr[1],
		GW_Ptr[0] }), 
	.SYNC({ GW_Ptr_Syn[3],
		GW_Ptr_Syn[2],
		GW_Ptr_Syn[1],
		GW_Ptr_Syn[0] }), 
	.test_se(test_se), 
	.FE_OFN5_M_Domain2_SYNC_RST(FE_OFN5_M_Domain2_SYNC_RST), 
	.TX_CLK_M__L3_N3(TX_CLK_M__L3_N3));
   FIFO_R_Addr_Size3_test_1 U2_FIFO_R (.R_CLK(I_R_CLK), 
	.R_RST(I_R_RST), 
	.R_INC(I_R_INC), 
	.GW_Ptr_Syn({ GW_Ptr_Syn[3],
		GW_Ptr_Syn[2],
		GW_Ptr_Syn[1],
		GW_Ptr_Syn[0] }), 
	.FIFO_Empty(FIFO_Empty), 
	.R_Addr({ R_Addr[2],
		R_Addr[1],
		R_Addr[0] }), 
	.GR_Ptr({ GR_Ptr[3],
		GR_Ptr[2],
		GR_Ptr[1],
		GR_Ptr[0] }), 
	.test_se(test_se), 
	.FE_OFN5_M_Domain2_SYNC_RST(FE_OFN5_M_Domain2_SYNC_RST), 
	.TX_CLK_M__L3_N3(TX_CLK_M__L3_N3));
   BIT_SYNC_2_00000004_test_1 U3_R2W_SYNC (.CLK(REF_CLK_M__L5_N4), 
	.RST(I_W_RST), 
	.ASYNC({ GR_Ptr[3],
		GR_Ptr[2],
		GR_Ptr[1],
		GR_Ptr[0] }), 
	.SYNC({ GR_Ptr_Syn[3],
		GR_Ptr_Syn[2],
		GR_Ptr_Syn[1],
		GR_Ptr_Syn[0] }), 
	.test_se(test_se));
   FIFO_MEM_Data_Width8_Addr_Size3_FIFO_Dipth8_test_1 U4_FIFO_MEM (.W_CLK(I_W_CLK), 
	.W_RST(I_W_RST), 
	.W_INC(I_W_INC), 
	.FIFO_Full(FIFO_Full), 
	.W_Addr({ W_Addr[2],
		W_Addr[1],
		W_Addr[0] }), 
	.W_Data({ I_Data[7],
		I_Data[6],
		I_Data[5],
		I_Data[4],
		I_Data[3],
		I_Data[2],
		I_Data[1],
		I_Data[0] }), 
	.R_Addr({ R_Addr[2],
		R_Addr[1],
		R_Addr[0] }), 
	.R_Data({ O_Data[7],
		O_Data[6],
		O_Data[5],
		O_Data[4],
		O_Data[3],
		O_Data[2],
		O_Data[1],
		O_Data[0] }), 
	.test_si2(test_si2), 
	.test_si1(GR_Ptr_Syn[3]), 
	.test_so2(test_so2), 
	.test_so1(test_so1), 
	.test_se(test_se), 
	.FE_OFN1_M_Domain1_SYNC_RST(FE_OFN1_M_Domain1_SYNC_RST), 
	.FE_OFN4_M_Domain1_SYNC_RST(FE_OFN4_M_Domain1_SYNC_RST), 
	.REF_CLK_M__L5_N1(REF_CLK_M__L5_N1), 
	.REF_CLK_M__L5_N4(REF_CLK_M__L5_N4), 
	.REF_CLK_M__L5_N5(REF_CLK_M__L5_N5), 
	.REF_CLK_M__L5_N6(REF_CLK_M__L5_N6), 
	.REF_CLK_M__L5_N7(REF_CLK_M__L5_N7));
endmodule

module PULSE_GEN_test_1 (
	clk, 
	rst, 
	lvl_sig, 
	pulse_sig, 
	test_si, 
	test_so, 
	test_se);
   input clk;
   input rst;
   input lvl_sig;
   output pulse_sig;
   input test_si;
   output test_so;
   input test_se;

   // Internal wires
   wire pls_flop;
   wire rcv_flop;

   assign test_so = rcv_flop ;

   SDFFRQX2M rcv_flop_reg (.SI(pls_flop), 
	.SE(test_se), 
	.RN(rst), 
	.Q(rcv_flop), 
	.D(lvl_sig), 
	.CK(clk));
   SDFFRQX2M pls_flop_reg (.SI(test_si), 
	.SE(test_se), 
	.RN(rst), 
	.Q(pls_flop), 
	.D(rcv_flop), 
	.CK(clk));
   NOR2BX2M U5 (.Y(pulse_sig), 
	.B(pls_flop), 
	.AN(rcv_flop));
endmodule

module RST_SYN_NUM_STAGES2_test_0 (
	RST, 
	CLK, 
	SYNC_RST, 
	test_si, 
	test_se);
   input RST;
   input CLK;
   output SYNC_RST;
   input test_si;
   input test_se;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire \sync_reg[0] ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   SDFFRQX2M \sync_reg_reg[1]  (.SI(\sync_reg[0] ), 
	.SE(test_se), 
	.RN(RST), 
	.Q(SYNC_RST), 
	.D(\sync_reg[0] ), 
	.CK(CLK));
   SDFFRQX2M \sync_reg_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.Q(\sync_reg[0] ), 
	.D(HTIE_LTIEHI_NET), 
	.CK(CLK));
endmodule

module RST_SYN_NUM_STAGES2_test_1 (
	RST, 
	CLK, 
	SYNC_RST, 
	test_si, 
	test_se);
   input RST;
   input CLK;
   output SYNC_RST;
   input test_si;
   input test_se;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire \sync_reg[0] ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   SDFFRQX2M \sync_reg_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.Q(\sync_reg[0] ), 
	.D(HTIE_LTIEHI_NET), 
	.CK(CLK));
   SDFFRQX1M \sync_reg_reg[1]  (.SI(\sync_reg[0] ), 
	.SE(test_se), 
	.RN(RST), 
	.Q(SYNC_RST), 
	.D(\sync_reg[0] ), 
	.CK(CLK));
endmodule

module DATA_SYNC_NUM_STAGES2_BUS_WIDTH8_test_1 (
	CLK, 
	RST, 
	unsync_bus, 
	bus_enable, 
	sync_bus, 
	enable_pulse_d, 
	test_si, 
	test_se, 
	REF_CLK_M__L5_N2, 
	REF_CLK_M__L5_N3);
   input CLK;
   input RST;
   input [7:0] unsync_bus;
   input bus_enable;
   output [7:0] sync_bus;
   output enable_pulse_d;
   input test_si;
   input test_se;
   input REF_CLK_M__L5_N2;
   input REF_CLK_M__L5_N3;

   // Internal wires
   wire Pulse_FF_Out;
   wire n1;
   wire n4;
   wire n6;
   wire n8;
   wire n10;
   wire n12;
   wire n14;
   wire n16;
   wire n18;
   wire n22;
   wire [1:0] en_sync_reg;

   SDFFRQX2M Pulse_FF_Out_reg (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.Q(Pulse_FF_Out), 
	.D(en_sync_reg[1]), 
	.CK(CLK));
   SDFFRQX2M \en_sync_reg_reg[1]  (.SI(en_sync_reg[0]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(en_sync_reg[1]), 
	.D(en_sync_reg[0]), 
	.CK(CLK));
   SDFFRQX2M \sync_bus_reg[3]  (.SI(sync_bus[2]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(sync_bus[3]), 
	.D(n10), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \sync_bus_reg[7]  (.SI(sync_bus[6]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(sync_bus[7]), 
	.D(n18), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \sync_bus_reg[4]  (.SI(sync_bus[3]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(sync_bus[4]), 
	.D(n12), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \sync_bus_reg[0]  (.SI(enable_pulse_d), 
	.SE(test_se), 
	.RN(RST), 
	.Q(sync_bus[0]), 
	.D(n4), 
	.CK(CLK));
   SDFFRQX2M \sync_bus_reg[2]  (.SI(sync_bus[1]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(sync_bus[2]), 
	.D(n8), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \sync_bus_reg[1]  (.SI(sync_bus[0]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(sync_bus[1]), 
	.D(n6), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \sync_bus_reg[6]  (.SI(sync_bus[5]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(sync_bus[6]), 
	.D(n16), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \sync_bus_reg[5]  (.SI(sync_bus[4]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(sync_bus[5]), 
	.D(n14), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M enable_pulse_d_reg (.SI(en_sync_reg[1]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(enable_pulse_d), 
	.D(n22), 
	.CK(CLK));
   SDFFRQX2M \en_sync_reg_reg[0]  (.SI(Pulse_FF_Out), 
	.SE(test_se), 
	.RN(RST), 
	.Q(en_sync_reg[0]), 
	.D(bus_enable), 
	.CK(CLK));
   INVX2M U3 (.Y(n22), 
	.A(n1));
   NAND2BX2M U4 (.Y(n1), 
	.B(en_sync_reg[1]), 
	.AN(Pulse_FF_Out));
   AO22X1M U5 (.Y(n4), 
	.B1(n1), 
	.B0(sync_bus[0]), 
	.A1(n22), 
	.A0(unsync_bus[0]));
   AO22X1M U6 (.Y(n6), 
	.B1(n1), 
	.B0(sync_bus[1]), 
	.A1(n22), 
	.A0(unsync_bus[1]));
   AO22X1M U7 (.Y(n8), 
	.B1(n1), 
	.B0(sync_bus[2]), 
	.A1(n22), 
	.A0(unsync_bus[2]));
   AO22X1M U8 (.Y(n10), 
	.B1(n1), 
	.B0(sync_bus[3]), 
	.A1(n22), 
	.A0(unsync_bus[3]));
   AO22X1M U9 (.Y(n12), 
	.B1(n1), 
	.B0(sync_bus[4]), 
	.A1(n22), 
	.A0(unsync_bus[4]));
   AO22X1M U10 (.Y(n14), 
	.B1(n1), 
	.B0(sync_bus[5]), 
	.A1(n22), 
	.A0(unsync_bus[5]));
   AO22X1M U11 (.Y(n16), 
	.B1(n1), 
	.B0(sync_bus[6]), 
	.A1(n22), 
	.A0(unsync_bus[6]));
   AO22X1M U12 (.Y(n18), 
	.B1(n1), 
	.B0(sync_bus[7]), 
	.A1(n22), 
	.A0(unsync_bus[7]));
endmodule

module CLK_GATE (
	CLK_EN, 
	CLK, 
	GATED_CLK);
   input CLK_EN;
   input CLK;
   output GATED_CLK;

   TLATNCAX12M U0_TLATNCAX12M (.ECK(GATED_CLK), 
	.E(CLK_EN), 
	.CK(CLK));
endmodule

module ALU_IN_Width8_DW_div_uns_0 (
	a, 
	b, 
	quotient, 
	remainder, 
	divide_by_0, 
	n144, 
	n151, 
	n152, 
	n149, 
	n150, 
	n160, 
	n143, 
	n159, 
	n158, 
	n157, 
	n156, 
	n155, 
	n148, 
	n147);
   input [7:0] a;
   input [7:0] b;
   output [7:0] quotient;
   output [7:0] remainder;
   output divide_by_0;
   input n144;
   input n151;
   input n152;
   input n149;
   input n150;
   input n160;
   input n143;
   input n159;
   input n158;
   input n157;
   input n156;
   input n155;
   input n148;
   input n147;

   // Internal wires
   wire \u_div/SumTmp[1][0] ;
   wire \u_div/SumTmp[1][1] ;
   wire \u_div/SumTmp[1][2] ;
   wire \u_div/SumTmp[1][3] ;
   wire \u_div/SumTmp[1][4] ;
   wire \u_div/SumTmp[1][5] ;
   wire \u_div/SumTmp[1][6] ;
   wire \u_div/SumTmp[2][0] ;
   wire \u_div/SumTmp[2][1] ;
   wire \u_div/SumTmp[2][2] ;
   wire \u_div/SumTmp[2][3] ;
   wire \u_div/SumTmp[2][4] ;
   wire \u_div/SumTmp[2][5] ;
   wire \u_div/SumTmp[3][0] ;
   wire \u_div/SumTmp[3][1] ;
   wire \u_div/SumTmp[3][2] ;
   wire \u_div/SumTmp[3][3] ;
   wire \u_div/SumTmp[3][4] ;
   wire \u_div/SumTmp[4][0] ;
   wire \u_div/SumTmp[4][1] ;
   wire \u_div/SumTmp[4][2] ;
   wire \u_div/SumTmp[4][3] ;
   wire \u_div/SumTmp[5][0] ;
   wire \u_div/SumTmp[5][1] ;
   wire \u_div/SumTmp[5][2] ;
   wire \u_div/SumTmp[6][0] ;
   wire \u_div/SumTmp[6][1] ;
   wire \u_div/SumTmp[7][0] ;
   wire \u_div/CryTmp[0][1] ;
   wire \u_div/CryTmp[0][2] ;
   wire \u_div/CryTmp[0][3] ;
   wire \u_div/CryTmp[0][4] ;
   wire \u_div/CryTmp[0][5] ;
   wire \u_div/CryTmp[0][6] ;
   wire \u_div/CryTmp[0][7] ;
   wire \u_div/CryTmp[1][1] ;
   wire \u_div/CryTmp[1][2] ;
   wire \u_div/CryTmp[1][3] ;
   wire \u_div/CryTmp[1][4] ;
   wire \u_div/CryTmp[1][5] ;
   wire \u_div/CryTmp[1][6] ;
   wire \u_div/CryTmp[1][7] ;
   wire \u_div/CryTmp[2][1] ;
   wire \u_div/CryTmp[2][2] ;
   wire \u_div/CryTmp[2][3] ;
   wire \u_div/CryTmp[2][4] ;
   wire \u_div/CryTmp[2][5] ;
   wire \u_div/CryTmp[2][6] ;
   wire \u_div/CryTmp[3][1] ;
   wire \u_div/CryTmp[3][2] ;
   wire \u_div/CryTmp[3][3] ;
   wire \u_div/CryTmp[3][4] ;
   wire \u_div/CryTmp[3][5] ;
   wire \u_div/CryTmp[4][1] ;
   wire \u_div/CryTmp[4][2] ;
   wire \u_div/CryTmp[4][3] ;
   wire \u_div/CryTmp[4][4] ;
   wire \u_div/CryTmp[5][1] ;
   wire \u_div/CryTmp[5][2] ;
   wire \u_div/CryTmp[5][3] ;
   wire \u_div/CryTmp[6][1] ;
   wire \u_div/CryTmp[6][2] ;
   wire \u_div/CryTmp[7][1] ;
   wire \u_div/PartRem[1][1] ;
   wire \u_div/PartRem[1][2] ;
   wire \u_div/PartRem[1][3] ;
   wire \u_div/PartRem[1][4] ;
   wire \u_div/PartRem[1][5] ;
   wire \u_div/PartRem[1][6] ;
   wire \u_div/PartRem[1][7] ;
   wire \u_div/PartRem[2][1] ;
   wire \u_div/PartRem[2][2] ;
   wire \u_div/PartRem[2][3] ;
   wire \u_div/PartRem[2][4] ;
   wire \u_div/PartRem[2][5] ;
   wire \u_div/PartRem[2][6] ;
   wire \u_div/PartRem[3][1] ;
   wire \u_div/PartRem[3][2] ;
   wire \u_div/PartRem[3][3] ;
   wire \u_div/PartRem[3][4] ;
   wire \u_div/PartRem[3][5] ;
   wire \u_div/PartRem[4][1] ;
   wire \u_div/PartRem[4][2] ;
   wire \u_div/PartRem[4][3] ;
   wire \u_div/PartRem[4][4] ;
   wire \u_div/PartRem[5][1] ;
   wire \u_div/PartRem[5][2] ;
   wire \u_div/PartRem[5][3] ;
   wire \u_div/PartRem[6][1] ;
   wire \u_div/PartRem[6][2] ;
   wire \u_div/PartRem[7][1] ;
   wire n1;
   wire n2;
   wire n3;
   wire n5;
   wire n7;
   wire n8;
   wire n9;
   wire n13;
   wire n14;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;

   ADDFX2M \u_div/u_fa_PartRem_0_2_5  (.S(\u_div/SumTmp[2][5] ), 
	.CO(\u_div/CryTmp[2][6] ), 
	.CI(\u_div/CryTmp[2][5] ), 
	.B(n13), 
	.A(\u_div/PartRem[3][5] ));
   ADDFX2M \u_div/u_fa_PartRem_0_4_3  (.S(\u_div/SumTmp[4][3] ), 
	.CO(\u_div/CryTmp[4][4] ), 
	.CI(\u_div/CryTmp[4][3] ), 
	.B(n151), 
	.A(\u_div/PartRem[5][3] ));
   ADDFX2M \u_div/u_fa_PartRem_0_5_2  (.S(\u_div/SumTmp[5][2] ), 
	.CO(\u_div/CryTmp[5][3] ), 
	.CI(\u_div/CryTmp[5][2] ), 
	.B(n16), 
	.A(\u_div/PartRem[6][2] ));
   ADDFX2M \u_div/u_fa_PartRem_0_6_1  (.S(\u_div/SumTmp[6][1] ), 
	.CO(\u_div/CryTmp[6][2] ), 
	.CI(\u_div/CryTmp[6][1] ), 
	.B(n17), 
	.A(\u_div/PartRem[7][1] ));
   ADDFX2M \u_div/u_fa_PartRem_0_3_4  (.S(\u_div/SumTmp[3][4] ), 
	.CO(\u_div/CryTmp[3][5] ), 
	.CI(\u_div/CryTmp[3][4] ), 
	.B(n14), 
	.A(\u_div/PartRem[4][4] ));
   ADDFX2M \u_div/u_fa_PartRem_0_0_6  (.CO(\u_div/CryTmp[0][7] ), 
	.CI(\u_div/CryTmp[0][6] ), 
	.B(n148), 
	.A(\u_div/PartRem[1][6] ));
   ADDFX2M \u_div/u_fa_PartRem_0_0_7  (.CO(quotient[0]), 
	.CI(\u_div/CryTmp[0][7] ), 
	.B(n147), 
	.A(\u_div/PartRem[1][7] ));
   ADDFX2M \u_div/u_fa_PartRem_0_1_1  (.S(\u_div/SumTmp[1][1] ), 
	.CO(\u_div/CryTmp[1][2] ), 
	.CI(\u_div/CryTmp[1][1] ), 
	.B(n17), 
	.A(\u_div/PartRem[2][1] ));
   ADDFX2M \u_div/u_fa_PartRem_0_2_1  (.S(\u_div/SumTmp[2][1] ), 
	.CO(\u_div/CryTmp[2][2] ), 
	.CI(\u_div/CryTmp[2][1] ), 
	.B(n17), 
	.A(\u_div/PartRem[3][1] ));
   ADDFX2M \u_div/u_fa_PartRem_0_3_1  (.S(\u_div/SumTmp[3][1] ), 
	.CO(\u_div/CryTmp[3][2] ), 
	.CI(\u_div/CryTmp[3][1] ), 
	.B(n17), 
	.A(\u_div/PartRem[4][1] ));
   ADDFX2M \u_div/u_fa_PartRem_0_4_1  (.S(\u_div/SumTmp[4][1] ), 
	.CO(\u_div/CryTmp[4][2] ), 
	.CI(\u_div/CryTmp[4][1] ), 
	.B(n17), 
	.A(\u_div/PartRem[5][1] ));
   ADDFX2M \u_div/u_fa_PartRem_0_5_1  (.S(\u_div/SumTmp[5][1] ), 
	.CO(\u_div/CryTmp[5][2] ), 
	.CI(\u_div/CryTmp[5][1] ), 
	.B(n17), 
	.A(\u_div/PartRem[6][1] ));
   ADDFX2M \u_div/u_fa_PartRem_0_0_3  (.CO(\u_div/CryTmp[0][4] ), 
	.CI(\u_div/CryTmp[0][3] ), 
	.B(n151), 
	.A(\u_div/PartRem[1][3] ));
   ADDFX2M \u_div/u_fa_PartRem_0_0_4  (.CO(\u_div/CryTmp[0][5] ), 
	.CI(\u_div/CryTmp[0][4] ), 
	.B(n14), 
	.A(\u_div/PartRem[1][4] ));
   ADDFX2M \u_div/u_fa_PartRem_0_0_5  (.CO(\u_div/CryTmp[0][6] ), 
	.CI(\u_div/CryTmp[0][5] ), 
	.B(n13), 
	.A(\u_div/PartRem[1][5] ));
   ADDFX2M \u_div/u_fa_PartRem_0_1_4  (.S(\u_div/SumTmp[1][4] ), 
	.CO(\u_div/CryTmp[1][5] ), 
	.CI(\u_div/CryTmp[1][4] ), 
	.B(n14), 
	.A(\u_div/PartRem[2][4] ));
   ADDFX2M \u_div/u_fa_PartRem_0_0_1  (.CO(\u_div/CryTmp[0][2] ), 
	.CI(\u_div/CryTmp[0][1] ), 
	.B(n17), 
	.A(\u_div/PartRem[1][1] ));
   ADDFX2M \u_div/u_fa_PartRem_0_0_2  (.CO(\u_div/CryTmp[0][3] ), 
	.CI(\u_div/CryTmp[0][2] ), 
	.B(n16), 
	.A(\u_div/PartRem[1][2] ));
   ADDFX2M \u_div/u_fa_PartRem_0_1_3  (.S(\u_div/SumTmp[1][3] ), 
	.CO(\u_div/CryTmp[1][4] ), 
	.CI(\u_div/CryTmp[1][3] ), 
	.B(n151), 
	.A(\u_div/PartRem[2][3] ));
   ADDFX2M \u_div/u_fa_PartRem_0_1_5  (.S(\u_div/SumTmp[1][5] ), 
	.CO(\u_div/CryTmp[1][6] ), 
	.CI(\u_div/CryTmp[1][5] ), 
	.B(n13), 
	.A(\u_div/PartRem[2][5] ));
   ADDFX2M \u_div/u_fa_PartRem_0_1_2  (.S(\u_div/SumTmp[1][2] ), 
	.CO(\u_div/CryTmp[1][3] ), 
	.CI(\u_div/CryTmp[1][2] ), 
	.B(n16), 
	.A(\u_div/PartRem[2][2] ));
   ADDFX2M \u_div/u_fa_PartRem_0_2_4  (.S(\u_div/SumTmp[2][4] ), 
	.CO(\u_div/CryTmp[2][5] ), 
	.CI(\u_div/CryTmp[2][4] ), 
	.B(n14), 
	.A(\u_div/PartRem[3][4] ));
   ADDFX2M \u_div/u_fa_PartRem_0_2_3  (.S(\u_div/SumTmp[2][3] ), 
	.CO(\u_div/CryTmp[2][4] ), 
	.CI(\u_div/CryTmp[2][3] ), 
	.B(n151), 
	.A(\u_div/PartRem[3][3] ));
   ADDFX2M \u_div/u_fa_PartRem_0_2_2  (.S(\u_div/SumTmp[2][2] ), 
	.CO(\u_div/CryTmp[2][3] ), 
	.CI(\u_div/CryTmp[2][2] ), 
	.B(n16), 
	.A(\u_div/PartRem[3][2] ));
   ADDFX2M \u_div/u_fa_PartRem_0_3_3  (.S(\u_div/SumTmp[3][3] ), 
	.CO(\u_div/CryTmp[3][4] ), 
	.CI(\u_div/CryTmp[3][3] ), 
	.B(n151), 
	.A(\u_div/PartRem[4][3] ));
   ADDFX2M \u_div/u_fa_PartRem_0_3_2  (.S(\u_div/SumTmp[3][2] ), 
	.CO(\u_div/CryTmp[3][3] ), 
	.CI(\u_div/CryTmp[3][2] ), 
	.B(n16), 
	.A(\u_div/PartRem[4][2] ));
   ADDFX2M \u_div/u_fa_PartRem_0_4_2  (.S(\u_div/SumTmp[4][2] ), 
	.CO(\u_div/CryTmp[4][3] ), 
	.CI(\u_div/CryTmp[4][2] ), 
	.B(n16), 
	.A(\u_div/PartRem[5][2] ));
   ADDFX2M \u_div/u_fa_PartRem_0_1_6  (.S(\u_div/SumTmp[1][6] ), 
	.CO(\u_div/CryTmp[1][7] ), 
	.CI(\u_div/CryTmp[1][6] ), 
	.B(n148), 
	.A(\u_div/PartRem[2][6] ));
   INVX2M U1 (.Y(n18), 
	.A(b[0]));
   XNOR2X2M U2 (.Y(\u_div/SumTmp[7][0] ), 
	.B(a[7]), 
	.A(n18));
   XNOR2X2M U3 (.Y(\u_div/SumTmp[6][0] ), 
	.B(a[6]), 
	.A(n18));
   XNOR2X2M U4 (.Y(\u_div/SumTmp[5][0] ), 
	.B(a[5]), 
	.A(n18));
   XNOR2X2M U5 (.Y(\u_div/SumTmp[4][0] ), 
	.B(a[4]), 
	.A(n18));
   XNOR2X2M U6 (.Y(\u_div/SumTmp[3][0] ), 
	.B(a[3]), 
	.A(n18));
   XNOR2X2M U7 (.Y(\u_div/SumTmp[2][0] ), 
	.B(a[2]), 
	.A(n18));
   XNOR2X2M U8 (.Y(\u_div/SumTmp[1][0] ), 
	.B(a[1]), 
	.A(n18));
   OR2X2M U9 (.Y(\u_div/CryTmp[7][1] ), 
	.B(a[7]), 
	.A(n18));
   INVX2M U10 (.Y(n17), 
	.A(b[1]));
   NAND2X2M U11 (.Y(\u_div/CryTmp[0][1] ), 
	.B(n160), 
	.A(n2));
   NAND2X2M U12 (.Y(\u_div/CryTmp[5][1] ), 
	.B(n3), 
	.A(n2));
   INVX2M U13 (.Y(n3), 
	.A(a[5]));
   INVX2M U14 (.Y(n2), 
	.A(n18));
   NAND2X2M U15 (.Y(\u_div/CryTmp[4][1] ), 
	.B(n5), 
	.A(n2));
   INVX2M U16 (.Y(n5), 
	.A(a[4]));
   NAND2X2M U18 (.Y(\u_div/CryTmp[3][1] ), 
	.B(n7), 
	.A(n2));
   INVX2M U19 (.Y(n7), 
	.A(a[3]));
   NAND2X2M U21 (.Y(\u_div/CryTmp[2][1] ), 
	.B(n8), 
	.A(n2));
   INVX2M U22 (.Y(n8), 
	.A(a[2]));
   NAND2X2M U23 (.Y(\u_div/CryTmp[1][1] ), 
	.B(n9), 
	.A(n2));
   INVX2M U24 (.Y(n9), 
	.A(a[1]));
   NAND2X2M U25 (.Y(\u_div/CryTmp[6][1] ), 
	.B(n1), 
	.A(n2));
   INVX2M U26 (.Y(n1), 
	.A(a[6]));
   INVX2M U30 (.Y(n16), 
	.A(b[2]));
   INVX2M U32 (.Y(n14), 
	.A(b[4]));
   INVX2M U33 (.Y(n13), 
	.A(b[5]));
   CLKMX2X2M U34 (.Y(\u_div/PartRem[1][7] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][6] ), 
	.A(\u_div/PartRem[2][6] ));
   CLKMX2X2M U35 (.Y(\u_div/PartRem[2][6] ), 
	.S0(quotient[2]), 
	.B(\u_div/SumTmp[2][5] ), 
	.A(\u_div/PartRem[3][5] ));
   CLKMX2X2M U36 (.Y(\u_div/PartRem[3][5] ), 
	.S0(quotient[3]), 
	.B(\u_div/SumTmp[3][4] ), 
	.A(\u_div/PartRem[4][4] ));
   CLKMX2X2M U37 (.Y(\u_div/PartRem[4][4] ), 
	.S0(quotient[4]), 
	.B(\u_div/SumTmp[4][3] ), 
	.A(\u_div/PartRem[5][3] ));
   CLKMX2X2M U38 (.Y(\u_div/PartRem[5][3] ), 
	.S0(quotient[5]), 
	.B(\u_div/SumTmp[5][2] ), 
	.A(\u_div/PartRem[6][2] ));
   CLKMX2X2M U39 (.Y(\u_div/PartRem[6][2] ), 
	.S0(quotient[6]), 
	.B(\u_div/SumTmp[6][1] ), 
	.A(\u_div/PartRem[7][1] ));
   CLKMX2X2M U40 (.Y(\u_div/PartRem[7][1] ), 
	.S0(quotient[7]), 
	.B(\u_div/SumTmp[7][0] ), 
	.A(a[7]));
   CLKMX2X2M U41 (.Y(\u_div/PartRem[1][6] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][5] ), 
	.A(\u_div/PartRem[2][5] ));
   CLKMX2X2M U42 (.Y(\u_div/PartRem[2][5] ), 
	.S0(quotient[2]), 
	.B(\u_div/SumTmp[2][4] ), 
	.A(\u_div/PartRem[3][4] ));
   CLKMX2X2M U43 (.Y(\u_div/PartRem[3][4] ), 
	.S0(quotient[3]), 
	.B(\u_div/SumTmp[3][3] ), 
	.A(\u_div/PartRem[4][3] ));
   CLKMX2X2M U44 (.Y(\u_div/PartRem[4][3] ), 
	.S0(quotient[4]), 
	.B(\u_div/SumTmp[4][2] ), 
	.A(\u_div/PartRem[5][2] ));
   CLKMX2X2M U45 (.Y(\u_div/PartRem[5][2] ), 
	.S0(quotient[5]), 
	.B(\u_div/SumTmp[5][1] ), 
	.A(\u_div/PartRem[6][1] ));
   CLKMX2X2M U46 (.Y(\u_div/PartRem[6][1] ), 
	.S0(quotient[6]), 
	.B(\u_div/SumTmp[6][0] ), 
	.A(a[6]));
   CLKMX2X2M U47 (.Y(\u_div/PartRem[1][5] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][4] ), 
	.A(\u_div/PartRem[2][4] ));
   CLKMX2X2M U48 (.Y(\u_div/PartRem[2][4] ), 
	.S0(quotient[2]), 
	.B(\u_div/SumTmp[2][3] ), 
	.A(\u_div/PartRem[3][3] ));
   CLKMX2X2M U49 (.Y(\u_div/PartRem[3][3] ), 
	.S0(quotient[3]), 
	.B(\u_div/SumTmp[3][2] ), 
	.A(\u_div/PartRem[4][2] ));
   CLKMX2X2M U50 (.Y(\u_div/PartRem[4][2] ), 
	.S0(quotient[4]), 
	.B(\u_div/SumTmp[4][1] ), 
	.A(\u_div/PartRem[5][1] ));
   CLKMX2X2M U51 (.Y(\u_div/PartRem[5][1] ), 
	.S0(quotient[5]), 
	.B(\u_div/SumTmp[5][0] ), 
	.A(a[5]));
   CLKMX2X2M U52 (.Y(\u_div/PartRem[1][4] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][3] ), 
	.A(\u_div/PartRem[2][3] ));
   CLKMX2X2M U53 (.Y(\u_div/PartRem[2][3] ), 
	.S0(quotient[2]), 
	.B(\u_div/SumTmp[2][2] ), 
	.A(\u_div/PartRem[3][2] ));
   CLKMX2X2M U54 (.Y(\u_div/PartRem[3][2] ), 
	.S0(quotient[3]), 
	.B(\u_div/SumTmp[3][1] ), 
	.A(\u_div/PartRem[4][1] ));
   CLKMX2X2M U55 (.Y(\u_div/PartRem[4][1] ), 
	.S0(quotient[4]), 
	.B(\u_div/SumTmp[4][0] ), 
	.A(a[4]));
   CLKMX2X2M U56 (.Y(\u_div/PartRem[1][3] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][2] ), 
	.A(\u_div/PartRem[2][2] ));
   CLKMX2X2M U57 (.Y(\u_div/PartRem[2][2] ), 
	.S0(quotient[2]), 
	.B(\u_div/SumTmp[2][1] ), 
	.A(\u_div/PartRem[3][1] ));
   CLKMX2X2M U58 (.Y(\u_div/PartRem[3][1] ), 
	.S0(quotient[3]), 
	.B(\u_div/SumTmp[3][0] ), 
	.A(a[3]));
   CLKMX2X2M U59 (.Y(\u_div/PartRem[1][2] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][1] ), 
	.A(\u_div/PartRem[2][1] ));
   CLKMX2X2M U60 (.Y(\u_div/PartRem[2][1] ), 
	.S0(quotient[2]), 
	.B(\u_div/SumTmp[2][0] ), 
	.A(a[2]));
   CLKMX2X2M U61 (.Y(\u_div/PartRem[1][1] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][0] ), 
	.A(a[1]));
   AND4X1M U62 (.Y(quotient[7]), 
	.D(n16), 
	.C(n17), 
	.B(n19), 
	.A(\u_div/CryTmp[7][1] ));
   AND3X1M U63 (.Y(quotient[6]), 
	.C(\u_div/CryTmp[6][2] ), 
	.B(n16), 
	.A(n19));
   AND2X1M U64 (.Y(quotient[5]), 
	.B(n19), 
	.A(\u_div/CryTmp[5][3] ));
   AND2X1M U65 (.Y(n19), 
	.B(n151), 
	.A(n20));
   AND2X1M U66 (.Y(quotient[4]), 
	.B(n20), 
	.A(\u_div/CryTmp[4][4] ));
   AND3X1M U67 (.Y(n20), 
	.C(n13), 
	.B(n14), 
	.A(n21));
   AND3X1M U68 (.Y(quotient[3]), 
	.C(\u_div/CryTmp[3][5] ), 
	.B(n13), 
	.A(n21));
   AND2X1M U69 (.Y(quotient[2]), 
	.B(n21), 
	.A(\u_div/CryTmp[2][6] ));
   NOR2X1M U70 (.Y(n21), 
	.B(b[7]), 
	.A(b[6]));
   AND2X1M U71 (.Y(quotient[1]), 
	.B(n147), 
	.A(\u_div/CryTmp[1][7] ));
endmodule

module ALU_IN_Width8_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO, 
	n144, 
	n151, 
	n152, 
	n149, 
	n150, 
	n160, 
	n148, 
	n147);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] DIFF;
   output CO;
   input n144;
   input n151;
   input n152;
   input n149;
   input n150;
   input n160;
   input n148;
   input n147;

   // Internal wires
   wire n4;
   wire n5;
   wire n7;
   wire n8;
   wire n9;
   wire [9:0] carry;

   ADDFX2M U2_5 (.S(DIFF[5]), 
	.CO(carry[6]), 
	.CI(carry[5]), 
	.B(n4), 
	.A(A[5]));
   ADDFX2M U2_4 (.S(DIFF[4]), 
	.CO(carry[5]), 
	.CI(carry[4]), 
	.B(n5), 
	.A(A[4]));
   ADDFX2M U2_3 (.S(DIFF[3]), 
	.CO(carry[4]), 
	.CI(carry[3]), 
	.B(n151), 
	.A(A[3]));
   ADDFX2M U2_2 (.S(DIFF[2]), 
	.CO(carry[3]), 
	.CI(carry[2]), 
	.B(n7), 
	.A(A[2]));
   ADDFX2M U2_7 (.S(DIFF[7]), 
	.CO(carry[8]), 
	.CI(carry[7]), 
	.B(n147), 
	.A(A[7]));
   ADDFX2M U2_1 (.S(DIFF[1]), 
	.CO(carry[2]), 
	.CI(carry[1]), 
	.B(n8), 
	.A(A[1]));
   ADDFX2M U2_6 (.S(DIFF[6]), 
	.CO(carry[7]), 
	.CI(carry[6]), 
	.B(n148), 
	.A(A[6]));
   XNOR2X2M U1 (.Y(DIFF[0]), 
	.B(A[0]), 
	.A(n9));
   INVX2M U3 (.Y(n8), 
	.A(B[1]));
   NAND2X2M U4 (.Y(carry[1]), 
	.B(n160), 
	.A(B[0]));
   INVX2M U7 (.Y(n9), 
	.A(B[0]));
   INVX2M U8 (.Y(n7), 
	.A(B[2]));
   INVX2M U10 (.Y(n5), 
	.A(B[4]));
   INVX2M U11 (.Y(n4), 
	.A(B[5]));
   CLKINVX1M U12 (.Y(DIFF[8]), 
	.A(carry[8]));
endmodule

module ALU_IN_Width8_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [8:1] carry;

   ADDFX2M U1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.CI(n1), 
	.B(B[1]), 
	.A(A[1]));
   ADDFX2M U1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.CI(carry[5]), 
	.B(B[5]), 
	.A(A[5]));
   ADDFX2M U1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.CI(carry[4]), 
	.B(B[4]), 
	.A(A[4]));
   ADDFX2M U1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.CI(carry[3]), 
	.B(B[3]), 
	.A(A[3]));
   ADDFX2M U1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.CI(carry[2]), 
	.B(B[2]), 
	.A(A[2]));
   ADDFX2M U1_7 (.S(SUM[7]), 
	.CO(SUM[8]), 
	.CI(carry[7]), 
	.B(B[7]), 
	.A(A[7]));
   ADDFX2M U1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.CI(carry[6]), 
	.B(B[6]), 
	.A(A[6]));
   AND2X2M U1 (.Y(n1), 
	.B(A[0]), 
	.A(B[0]));
   CLKXOR2X2M U2 (.Y(SUM[0]), 
	.B(A[0]), 
	.A(B[0]));
endmodule

module ALU_IN_Width8_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [13:0] A;
   input [13:0] B;
   input CI;
   output [13:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;

   AOI21BX2M U2 (.Y(n1), 
	.B0N(n19), 
	.A1(A[12]), 
	.A0(n18));
   NAND2X2M U3 (.Y(n15), 
	.B(B[7]), 
	.A(A[7]));
   XNOR2X2M U4 (.Y(SUM[7]), 
	.B(n8), 
	.A(A[7]));
   INVX2M U5 (.Y(n8), 
	.A(B[7]));
   XNOR2X2M U6 (.Y(SUM[13]), 
	.B(n1), 
	.A(B[13]));
   INVX2M U7 (.Y(n9), 
	.A(A[6]));
   INVX2M U8 (.Y(SUM[6]), 
	.A(n9));
   BUFX2M U9 (.Y(SUM[0]), 
	.A(A[0]));
   BUFX2M U10 (.Y(SUM[1]), 
	.A(A[1]));
   BUFX2M U11 (.Y(SUM[2]), 
	.A(A[2]));
   BUFX2M U12 (.Y(SUM[3]), 
	.A(A[3]));
   BUFX2M U13 (.Y(SUM[4]), 
	.A(A[4]));
   BUFX2M U14 (.Y(SUM[5]), 
	.A(A[5]));
   XNOR2X1M U15 (.Y(SUM[9]), 
	.B(n11), 
	.A(n10));
   NOR2X1M U16 (.Y(n11), 
	.B(n13), 
	.A(n12));
   CLKXOR2X2M U17 (.Y(SUM[8]), 
	.B(n15), 
	.A(n14));
   NAND2BX1M U18 (.Y(n14), 
	.B(n17), 
	.AN(n16));
   OAI21X1M U19 (.Y(n19), 
	.B0(B[12]), 
	.A1(n18), 
	.A0(A[12]));
   XOR3XLM U20 (.Y(SUM[12]), 
	.C(n18), 
	.B(A[12]), 
	.A(B[12]));
   OAI21BX1M U21 (.Y(n18), 
	.B0N(n22), 
	.A1(n21), 
	.A0(n20));
   XNOR2X1M U22 (.Y(SUM[11]), 
	.B(n23), 
	.A(n21));
   NOR2X1M U23 (.Y(n23), 
	.B(n20), 
	.A(n22));
   NOR2X1M U24 (.Y(n20), 
	.B(A[11]), 
	.A(B[11]));
   AND2X1M U25 (.Y(n22), 
	.B(A[11]), 
	.A(B[11]));
   OA21X1M U26 (.Y(n21), 
	.B0(n26), 
	.A1(n25), 
	.A0(n24));
   CLKXOR2X2M U27 (.Y(SUM[10]), 
	.B(n25), 
	.A(n27));
   AOI2BB1X1M U28 (.Y(n25), 
	.B0(n12), 
	.A1N(n13), 
	.A0N(n10));
   AND2X1M U29 (.Y(n12), 
	.B(A[9]), 
	.A(B[9]));
   NOR2X1M U30 (.Y(n13), 
	.B(A[9]), 
	.A(B[9]));
   OA21X1M U31 (.Y(n10), 
	.B0(n17), 
	.A1(n16), 
	.A0(n15));
   CLKNAND2X2M U32 (.Y(n17), 
	.B(A[8]), 
	.A(B[8]));
   NOR2X1M U33 (.Y(n16), 
	.B(A[8]), 
	.A(B[8]));
   NAND2BX1M U34 (.Y(n27), 
	.B(n26), 
	.AN(n24));
   CLKNAND2X2M U35 (.Y(n26), 
	.B(A[10]), 
	.A(B[10]));
   NOR2X1M U36 (.Y(n24), 
	.B(A[10]), 
	.A(B[10]));
endmodule

module ALU_IN_Width8_DW02_mult_0 (
	A, 
	B, 
	TC, 
	PRODUCT, 
	n144, 
	n151, 
	n152, 
	n149, 
	n150, 
	n160, 
	n143, 
	n159, 
	n158, 
	n157, 
	n156, 
	n155, 
	n154, 
	n148, 
	n147);
   input [7:0] A;
   input [7:0] B;
   input TC;
   output [15:0] PRODUCT;
   input n144;
   input n151;
   input n152;
   input n149;
   input n150;
   input n160;
   input n143;
   input n159;
   input n158;
   input n157;
   input n156;
   input n155;
   input n154;
   input n148;
   input n147;

   // Internal wires
   wire \ab[7][7] ;
   wire \ab[7][6] ;
   wire \ab[7][5] ;
   wire \ab[7][4] ;
   wire \ab[7][3] ;
   wire \ab[7][2] ;
   wire \ab[7][1] ;
   wire \ab[7][0] ;
   wire \ab[6][7] ;
   wire \ab[6][6] ;
   wire \ab[6][5] ;
   wire \ab[6][4] ;
   wire \ab[6][3] ;
   wire \ab[6][2] ;
   wire \ab[6][1] ;
   wire \ab[6][0] ;
   wire \ab[5][7] ;
   wire \ab[5][6] ;
   wire \ab[5][5] ;
   wire \ab[5][4] ;
   wire \ab[5][3] ;
   wire \ab[5][2] ;
   wire \ab[5][1] ;
   wire \ab[5][0] ;
   wire \ab[4][7] ;
   wire \ab[4][6] ;
   wire \ab[4][5] ;
   wire \ab[4][4] ;
   wire \ab[4][3] ;
   wire \ab[4][2] ;
   wire \ab[4][1] ;
   wire \ab[4][0] ;
   wire \ab[3][7] ;
   wire \ab[3][6] ;
   wire \ab[3][5] ;
   wire \ab[3][4] ;
   wire \ab[3][3] ;
   wire \ab[3][2] ;
   wire \ab[3][1] ;
   wire \ab[3][0] ;
   wire \ab[2][7] ;
   wire \ab[2][6] ;
   wire \ab[2][5] ;
   wire \ab[2][4] ;
   wire \ab[2][3] ;
   wire \ab[2][2] ;
   wire \ab[2][1] ;
   wire \ab[2][0] ;
   wire \ab[1][7] ;
   wire \ab[1][6] ;
   wire \ab[1][5] ;
   wire \ab[1][4] ;
   wire \ab[1][3] ;
   wire \ab[1][2] ;
   wire \ab[1][1] ;
   wire \ab[1][0] ;
   wire \ab[0][7] ;
   wire \ab[0][6] ;
   wire \ab[0][5] ;
   wire \ab[0][4] ;
   wire \ab[0][3] ;
   wire \ab[0][2] ;
   wire \ab[0][1] ;
   wire \CARRYB[7][6] ;
   wire \CARRYB[7][5] ;
   wire \CARRYB[7][4] ;
   wire \CARRYB[7][3] ;
   wire \CARRYB[7][2] ;
   wire \CARRYB[7][1] ;
   wire \CARRYB[7][0] ;
   wire \CARRYB[6][6] ;
   wire \CARRYB[6][5] ;
   wire \CARRYB[6][4] ;
   wire \CARRYB[6][3] ;
   wire \CARRYB[6][2] ;
   wire \CARRYB[6][1] ;
   wire \CARRYB[6][0] ;
   wire \CARRYB[5][6] ;
   wire \CARRYB[5][5] ;
   wire \CARRYB[5][4] ;
   wire \CARRYB[5][3] ;
   wire \CARRYB[5][2] ;
   wire \CARRYB[5][1] ;
   wire \CARRYB[5][0] ;
   wire \CARRYB[4][6] ;
   wire \CARRYB[4][5] ;
   wire \CARRYB[4][4] ;
   wire \CARRYB[4][3] ;
   wire \CARRYB[4][2] ;
   wire \CARRYB[4][1] ;
   wire \CARRYB[4][0] ;
   wire \CARRYB[3][6] ;
   wire \CARRYB[3][5] ;
   wire \CARRYB[3][4] ;
   wire \CARRYB[3][3] ;
   wire \CARRYB[3][2] ;
   wire \CARRYB[3][1] ;
   wire \CARRYB[3][0] ;
   wire \CARRYB[2][6] ;
   wire \CARRYB[2][5] ;
   wire \CARRYB[2][4] ;
   wire \CARRYB[2][3] ;
   wire \CARRYB[2][2] ;
   wire \CARRYB[2][1] ;
   wire \CARRYB[2][0] ;
   wire \SUMB[7][6] ;
   wire \SUMB[7][5] ;
   wire \SUMB[7][4] ;
   wire \SUMB[7][3] ;
   wire \SUMB[7][2] ;
   wire \SUMB[7][1] ;
   wire \SUMB[7][0] ;
   wire \SUMB[6][6] ;
   wire \SUMB[6][5] ;
   wire \SUMB[6][4] ;
   wire \SUMB[6][3] ;
   wire \SUMB[6][2] ;
   wire \SUMB[6][1] ;
   wire \SUMB[5][6] ;
   wire \SUMB[5][5] ;
   wire \SUMB[5][4] ;
   wire \SUMB[5][3] ;
   wire \SUMB[5][2] ;
   wire \SUMB[5][1] ;
   wire \SUMB[4][6] ;
   wire \SUMB[4][5] ;
   wire \SUMB[4][4] ;
   wire \SUMB[4][3] ;
   wire \SUMB[4][2] ;
   wire \SUMB[4][1] ;
   wire \SUMB[3][6] ;
   wire \SUMB[3][5] ;
   wire \SUMB[3][4] ;
   wire \SUMB[3][3] ;
   wire \SUMB[3][2] ;
   wire \SUMB[3][1] ;
   wire \SUMB[2][6] ;
   wire \SUMB[2][5] ;
   wire \SUMB[2][4] ;
   wire \SUMB[2][3] ;
   wire \SUMB[2][2] ;
   wire \SUMB[2][1] ;
   wire \SUMB[1][6] ;
   wire \SUMB[1][5] ;
   wire \SUMB[1][4] ;
   wire \SUMB[1][3] ;
   wire \SUMB[1][2] ;
   wire \SUMB[1][1] ;
   wire \A1[12] ;
   wire \A1[11] ;
   wire \A1[10] ;
   wire \A1[9] ;
   wire \A1[8] ;
   wire \A1[7] ;
   wire \A1[6] ;
   wire \A1[4] ;
   wire \A1[3] ;
   wire \A1[2] ;
   wire \A1[1] ;
   wire \A1[0] ;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n26;
   wire n27;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;

   ADDFX2M S1_6_0 (.S(\A1[4] ), 
	.CO(\CARRYB[6][0] ), 
	.CI(\SUMB[5][1] ), 
	.B(\CARRYB[5][0] ), 
	.A(\ab[6][0] ));
   ADDFX2M S1_5_0 (.S(\A1[3] ), 
	.CO(\CARRYB[5][0] ), 
	.CI(\SUMB[4][1] ), 
	.B(\CARRYB[4][0] ), 
	.A(\ab[5][0] ));
   ADDFX2M S1_4_0 (.S(\A1[2] ), 
	.CO(\CARRYB[4][0] ), 
	.CI(\SUMB[3][1] ), 
	.B(\CARRYB[3][0] ), 
	.A(\ab[4][0] ));
   ADDFX2M S1_3_0 (.S(\A1[1] ), 
	.CO(\CARRYB[3][0] ), 
	.CI(\SUMB[2][1] ), 
	.B(\CARRYB[2][0] ), 
	.A(\ab[3][0] ));
   ADDFX2M S2_6_5 (.S(\SUMB[6][5] ), 
	.CO(\CARRYB[6][5] ), 
	.CI(\SUMB[5][6] ), 
	.B(\CARRYB[5][5] ), 
	.A(\ab[6][5] ));
   ADDFX2M S2_6_4 (.S(\SUMB[6][4] ), 
	.CO(\CARRYB[6][4] ), 
	.CI(\SUMB[5][5] ), 
	.B(\CARRYB[5][4] ), 
	.A(\ab[6][4] ));
   ADDFX2M S2_5_5 (.S(\SUMB[5][5] ), 
	.CO(\CARRYB[5][5] ), 
	.CI(\SUMB[4][6] ), 
	.B(\CARRYB[4][5] ), 
	.A(\ab[5][5] ));
   ADDFX2M S2_6_3 (.S(\SUMB[6][3] ), 
	.CO(\CARRYB[6][3] ), 
	.CI(\SUMB[5][4] ), 
	.B(\CARRYB[5][3] ), 
	.A(\ab[6][3] ));
   ADDFX2M S2_5_4 (.S(\SUMB[5][4] ), 
	.CO(\CARRYB[5][4] ), 
	.CI(\SUMB[4][5] ), 
	.B(\CARRYB[4][4] ), 
	.A(\ab[5][4] ));
   ADDFX2M S2_6_2 (.S(\SUMB[6][2] ), 
	.CO(\CARRYB[6][2] ), 
	.CI(\SUMB[5][3] ), 
	.B(\CARRYB[5][2] ), 
	.A(\ab[6][2] ));
   ADDFX2M S2_4_5 (.S(\SUMB[4][5] ), 
	.CO(\CARRYB[4][5] ), 
	.CI(\SUMB[3][6] ), 
	.B(\CARRYB[3][5] ), 
	.A(\ab[4][5] ));
   ADDFX2M S2_5_2 (.S(\SUMB[5][2] ), 
	.CO(\CARRYB[5][2] ), 
	.CI(\SUMB[4][3] ), 
	.B(\CARRYB[4][2] ), 
	.A(\ab[5][2] ));
   ADDFX2M S2_5_3 (.S(\SUMB[5][3] ), 
	.CO(\CARRYB[5][3] ), 
	.CI(\SUMB[4][4] ), 
	.B(\CARRYB[4][3] ), 
	.A(\ab[5][3] ));
   ADDFX2M S2_4_2 (.S(\SUMB[4][2] ), 
	.CO(\CARRYB[4][2] ), 
	.CI(\SUMB[3][3] ), 
	.B(\CARRYB[3][2] ), 
	.A(\ab[4][2] ));
   ADDFX2M S2_4_3 (.S(\SUMB[4][3] ), 
	.CO(\CARRYB[4][3] ), 
	.CI(\SUMB[3][4] ), 
	.B(\CARRYB[3][3] ), 
	.A(\ab[4][3] ));
   ADDFX2M S2_4_4 (.S(\SUMB[4][4] ), 
	.CO(\CARRYB[4][4] ), 
	.CI(\SUMB[3][5] ), 
	.B(\CARRYB[3][4] ), 
	.A(\ab[4][4] ));
   ADDFX2M S2_3_2 (.S(\SUMB[3][2] ), 
	.CO(\CARRYB[3][2] ), 
	.CI(\SUMB[2][3] ), 
	.B(\CARRYB[2][2] ), 
	.A(\ab[3][2] ));
   ADDFX2M S2_3_3 (.S(\SUMB[3][3] ), 
	.CO(\CARRYB[3][3] ), 
	.CI(\SUMB[2][4] ), 
	.B(\CARRYB[2][3] ), 
	.A(\ab[3][3] ));
   ADDFX2M S2_3_4 (.S(\SUMB[3][4] ), 
	.CO(\CARRYB[3][4] ), 
	.CI(\SUMB[2][5] ), 
	.B(\CARRYB[2][4] ), 
	.A(\ab[3][4] ));
   ADDFX2M S2_3_5 (.S(\SUMB[3][5] ), 
	.CO(\CARRYB[3][5] ), 
	.CI(\SUMB[2][6] ), 
	.B(\CARRYB[2][5] ), 
	.A(\ab[3][5] ));
   ADDFX2M S1_2_0 (.S(\A1[0] ), 
	.CO(\CARRYB[2][0] ), 
	.CI(\SUMB[1][1] ), 
	.B(n9), 
	.A(\ab[2][0] ));
   ADDFX2M S2_2_2 (.S(\SUMB[2][2] ), 
	.CO(\CARRYB[2][2] ), 
	.CI(\SUMB[1][3] ), 
	.B(n8), 
	.A(\ab[2][2] ));
   ADDFX2M S2_2_3 (.S(\SUMB[2][3] ), 
	.CO(\CARRYB[2][3] ), 
	.CI(\SUMB[1][4] ), 
	.B(n7), 
	.A(\ab[2][3] ));
   ADDFX2M S2_2_4 (.S(\SUMB[2][4] ), 
	.CO(\CARRYB[2][4] ), 
	.CI(\SUMB[1][5] ), 
	.B(n6), 
	.A(\ab[2][4] ));
   ADDFX2M S2_2_5 (.S(\SUMB[2][5] ), 
	.CO(\CARRYB[2][5] ), 
	.CI(\SUMB[1][6] ), 
	.B(n5), 
	.A(\ab[2][5] ));
   ADDFX2M S4_0 (.S(\SUMB[7][0] ), 
	.CO(\CARRYB[7][0] ), 
	.CI(\SUMB[6][1] ), 
	.B(\CARRYB[6][0] ), 
	.A(\ab[7][0] ));
   ADDFX2M S4_5 (.S(\SUMB[7][5] ), 
	.CO(\CARRYB[7][5] ), 
	.CI(\SUMB[6][6] ), 
	.B(\CARRYB[6][5] ), 
	.A(\ab[7][5] ));
   ADDFX2M S4_4 (.S(\SUMB[7][4] ), 
	.CO(\CARRYB[7][4] ), 
	.CI(\SUMB[6][5] ), 
	.B(\CARRYB[6][4] ), 
	.A(\ab[7][4] ));
   ADDFX2M S4_3 (.S(\SUMB[7][3] ), 
	.CO(\CARRYB[7][3] ), 
	.CI(\SUMB[6][4] ), 
	.B(\CARRYB[6][3] ), 
	.A(\ab[7][3] ));
   ADDFX2M S4_2 (.S(\SUMB[7][2] ), 
	.CO(\CARRYB[7][2] ), 
	.CI(\SUMB[6][3] ), 
	.B(\CARRYB[6][2] ), 
	.A(\ab[7][2] ));
   ADDFX2M S2_6_1 (.S(\SUMB[6][1] ), 
	.CO(\CARRYB[6][1] ), 
	.CI(\SUMB[5][2] ), 
	.B(\CARRYB[5][1] ), 
	.A(\ab[6][1] ));
   ADDFX2M S2_5_1 (.S(\SUMB[5][1] ), 
	.CO(\CARRYB[5][1] ), 
	.CI(\SUMB[4][2] ), 
	.B(\CARRYB[4][1] ), 
	.A(\ab[5][1] ));
   ADDFX2M S2_4_1 (.S(\SUMB[4][1] ), 
	.CO(\CARRYB[4][1] ), 
	.CI(\SUMB[3][2] ), 
	.B(\CARRYB[3][1] ), 
	.A(\ab[4][1] ));
   ADDFX2M S2_3_1 (.S(\SUMB[3][1] ), 
	.CO(\CARRYB[3][1] ), 
	.CI(\SUMB[2][2] ), 
	.B(\CARRYB[2][1] ), 
	.A(\ab[3][1] ));
   ADDFX2M S3_6_6 (.S(\SUMB[6][6] ), 
	.CO(\CARRYB[6][6] ), 
	.CI(\ab[5][7] ), 
	.B(\CARRYB[5][6] ), 
	.A(\ab[6][6] ));
   ADDFX2M S3_5_6 (.S(\SUMB[5][6] ), 
	.CO(\CARRYB[5][6] ), 
	.CI(\ab[4][7] ), 
	.B(\CARRYB[4][6] ), 
	.A(\ab[5][6] ));
   ADDFX2M S3_4_6 (.S(\SUMB[4][6] ), 
	.CO(\CARRYB[4][6] ), 
	.CI(\ab[3][7] ), 
	.B(\CARRYB[3][6] ), 
	.A(\ab[4][6] ));
   ADDFX2M S3_3_6 (.S(\SUMB[3][6] ), 
	.CO(\CARRYB[3][6] ), 
	.CI(\ab[2][7] ), 
	.B(\CARRYB[2][6] ), 
	.A(\ab[3][6] ));
   ADDFX2M S3_2_6 (.S(\SUMB[2][6] ), 
	.CO(\CARRYB[2][6] ), 
	.CI(\ab[1][7] ), 
	.B(n4), 
	.A(\ab[2][6] ));
   ADDFX2M S2_2_1 (.S(\SUMB[2][1] ), 
	.CO(\CARRYB[2][1] ), 
	.CI(\SUMB[1][2] ), 
	.B(n3), 
	.A(\ab[2][1] ));
   ADDFX2M S5_6 (.S(\SUMB[7][6] ), 
	.CO(\CARRYB[7][6] ), 
	.CI(\ab[6][7] ), 
	.B(\CARRYB[6][6] ), 
	.A(\ab[7][6] ));
   ADDFX2M S4_1 (.S(\SUMB[7][1] ), 
	.CO(\CARRYB[7][1] ), 
	.CI(\SUMB[6][2] ), 
	.B(\CARRYB[6][1] ), 
	.A(\ab[7][1] ));
   AND2X2M U2 (.Y(n3), 
	.B(\ab[1][1] ), 
	.A(\ab[0][2] ));
   AND2X2M U3 (.Y(n4), 
	.B(\ab[1][6] ), 
	.A(\ab[0][7] ));
   AND2X2M U4 (.Y(n5), 
	.B(\ab[1][5] ), 
	.A(\ab[0][6] ));
   AND2X2M U5 (.Y(n6), 
	.B(\ab[1][4] ), 
	.A(\ab[0][5] ));
   AND2X2M U6 (.Y(n7), 
	.B(\ab[1][3] ), 
	.A(\ab[0][4] ));
   AND2X2M U7 (.Y(n8), 
	.B(\ab[1][2] ), 
	.A(\ab[0][3] ));
   AND2X2M U8 (.Y(n9), 
	.B(\ab[1][0] ), 
	.A(\ab[0][1] ));
   AND2X2M U9 (.Y(n10), 
	.B(\ab[7][7] ), 
	.A(\CARRYB[7][6] ));
   CLKXOR2X2M U10 (.Y(\A1[12] ), 
	.B(\ab[7][7] ), 
	.A(\CARRYB[7][6] ));
   INVX2M U11 (.Y(n23), 
	.A(\ab[0][7] ));
   INVX2M U12 (.Y(n22), 
	.A(\ab[0][6] ));
   CLKXOR2X2M U13 (.Y(\A1[7] ), 
	.B(\SUMB[7][2] ), 
	.A(\CARRYB[7][1] ));
   CLKXOR2X2M U14 (.Y(PRODUCT[1]), 
	.B(\ab[0][1] ), 
	.A(\ab[1][0] ));
   CLKXOR2X2M U15 (.Y(\A1[8] ), 
	.B(\SUMB[7][3] ), 
	.A(\CARRYB[7][2] ));
   CLKXOR2X2M U16 (.Y(\A1[10] ), 
	.B(\SUMB[7][5] ), 
	.A(\CARRYB[7][4] ));
   CLKXOR2X2M U17 (.Y(\A1[9] ), 
	.B(\SUMB[7][4] ), 
	.A(\CARRYB[7][3] ));
   CLKXOR2X2M U18 (.Y(\A1[11] ), 
	.B(\SUMB[7][6] ), 
	.A(\CARRYB[7][5] ));
   INVX2M U19 (.Y(n21), 
	.A(\ab[0][5] ));
   INVX2M U20 (.Y(n20), 
	.A(\ab[0][4] ));
   INVX2M U21 (.Y(n19), 
	.A(\ab[0][3] ));
   INVX2M U22 (.Y(n18), 
	.A(\ab[0][2] ));
   XNOR2X2M U23 (.Y(\SUMB[1][2] ), 
	.B(n19), 
	.A(\ab[1][2] ));
   XNOR2X2M U24 (.Y(\A1[6] ), 
	.B(n17), 
	.A(\CARRYB[7][0] ));
   INVX2M U25 (.Y(n17), 
	.A(\SUMB[7][1] ));
   AND2X2M U26 (.Y(n11), 
	.B(\SUMB[7][1] ), 
	.A(\CARRYB[7][0] ));
   AND2X2M U27 (.Y(n12), 
	.B(\SUMB[7][2] ), 
	.A(\CARRYB[7][1] ));
   AND2X2M U28 (.Y(n13), 
	.B(\SUMB[7][4] ), 
	.A(\CARRYB[7][3] ));
   AND2X2M U29 (.Y(n14), 
	.B(\SUMB[7][6] ), 
	.A(\CARRYB[7][5] ));
   AND2X2M U30 (.Y(n15), 
	.B(\SUMB[7][3] ), 
	.A(\CARRYB[7][2] ));
   AND2X2M U31 (.Y(n16), 
	.B(\SUMB[7][5] ), 
	.A(\CARRYB[7][4] ));
   XNOR2X2M U32 (.Y(\SUMB[1][6] ), 
	.B(n23), 
	.A(\ab[1][6] ));
   XNOR2X2M U33 (.Y(\SUMB[1][5] ), 
	.B(n22), 
	.A(\ab[1][5] ));
   XNOR2X2M U34 (.Y(\SUMB[1][4] ), 
	.B(n21), 
	.A(\ab[1][4] ));
   XNOR2X2M U35 (.Y(\SUMB[1][3] ), 
	.B(n20), 
	.A(\ab[1][3] ));
   XNOR2X2M U36 (.Y(\SUMB[1][1] ), 
	.B(n18), 
	.A(\ab[1][1] ));
   INVX2M U37 (.Y(n33), 
	.A(A[6]));
   INVX2M U38 (.Y(n32), 
	.A(A[7]));
   INVX2M U39 (.Y(n38), 
	.A(A[1]));
   INVX2M U41 (.Y(n37), 
	.A(A[2]));
   INVX2M U42 (.Y(n36), 
	.A(A[3]));
   INVX2M U44 (.Y(n34), 
	.A(A[5]));
   INVX2M U45 (.Y(n35), 
	.A(A[4]));
   INVX2M U47 (.Y(n30), 
	.A(B[1]));
   INVX2M U48 (.Y(n31), 
	.A(B[0]));
   INVX2M U50 (.Y(n29), 
	.A(B[2]));
   INVX2M U51 (.Y(n26), 
	.A(B[5]));
   INVX2M U52 (.Y(n27), 
	.A(B[4]));
   NOR2X1M U54 (.Y(\ab[7][7] ), 
	.B(n147), 
	.A(n32));
   NOR2X1M U55 (.Y(\ab[7][6] ), 
	.B(n148), 
	.A(n32));
   NOR2X1M U56 (.Y(\ab[7][5] ), 
	.B(n26), 
	.A(n32));
   NOR2X1M U57 (.Y(\ab[7][4] ), 
	.B(n27), 
	.A(n32));
   NOR2X1M U58 (.Y(\ab[7][3] ), 
	.B(n151), 
	.A(n32));
   NOR2X1M U59 (.Y(\ab[7][2] ), 
	.B(n29), 
	.A(n32));
   NOR2X1M U60 (.Y(\ab[7][1] ), 
	.B(n30), 
	.A(n32));
   NOR2X1M U61 (.Y(\ab[7][0] ), 
	.B(n31), 
	.A(n32));
   NOR2X1M U62 (.Y(\ab[6][7] ), 
	.B(n33), 
	.A(n147));
   NOR2X1M U63 (.Y(\ab[6][6] ), 
	.B(n33), 
	.A(n148));
   NOR2X1M U64 (.Y(\ab[6][5] ), 
	.B(n33), 
	.A(n26));
   NOR2X1M U65 (.Y(\ab[6][4] ), 
	.B(n33), 
	.A(n27));
   NOR2X1M U66 (.Y(\ab[6][3] ), 
	.B(n33), 
	.A(n151));
   NOR2X1M U67 (.Y(\ab[6][2] ), 
	.B(n33), 
	.A(n29));
   NOR2X1M U68 (.Y(\ab[6][1] ), 
	.B(n33), 
	.A(n30));
   NOR2X1M U69 (.Y(\ab[6][0] ), 
	.B(n33), 
	.A(n31));
   NOR2X1M U70 (.Y(\ab[5][7] ), 
	.B(n34), 
	.A(n147));
   NOR2X1M U71 (.Y(\ab[5][6] ), 
	.B(n34), 
	.A(n148));
   NOR2X1M U72 (.Y(\ab[5][5] ), 
	.B(n34), 
	.A(n26));
   NOR2X1M U73 (.Y(\ab[5][4] ), 
	.B(n34), 
	.A(n27));
   NOR2X1M U74 (.Y(\ab[5][3] ), 
	.B(n34), 
	.A(n151));
   NOR2X1M U75 (.Y(\ab[5][2] ), 
	.B(n34), 
	.A(n29));
   NOR2X1M U76 (.Y(\ab[5][1] ), 
	.B(n34), 
	.A(n30));
   NOR2X1M U77 (.Y(\ab[5][0] ), 
	.B(n34), 
	.A(n31));
   NOR2X1M U78 (.Y(\ab[4][7] ), 
	.B(n35), 
	.A(n147));
   NOR2X1M U79 (.Y(\ab[4][6] ), 
	.B(n35), 
	.A(n148));
   NOR2X1M U80 (.Y(\ab[4][5] ), 
	.B(n35), 
	.A(n26));
   NOR2X1M U81 (.Y(\ab[4][4] ), 
	.B(n35), 
	.A(n27));
   NOR2X1M U82 (.Y(\ab[4][3] ), 
	.B(n35), 
	.A(n151));
   NOR2X1M U83 (.Y(\ab[4][2] ), 
	.B(n35), 
	.A(n29));
   NOR2X1M U84 (.Y(\ab[4][1] ), 
	.B(n35), 
	.A(n30));
   NOR2X1M U85 (.Y(\ab[4][0] ), 
	.B(n35), 
	.A(n31));
   NOR2X1M U86 (.Y(\ab[3][7] ), 
	.B(n36), 
	.A(n147));
   NOR2X1M U87 (.Y(\ab[3][6] ), 
	.B(n36), 
	.A(n148));
   NOR2X1M U88 (.Y(\ab[3][5] ), 
	.B(n36), 
	.A(n26));
   NOR2X1M U89 (.Y(\ab[3][4] ), 
	.B(n36), 
	.A(n27));
   NOR2X1M U90 (.Y(\ab[3][3] ), 
	.B(n36), 
	.A(n151));
   NOR2X1M U91 (.Y(\ab[3][2] ), 
	.B(n36), 
	.A(n29));
   NOR2X1M U92 (.Y(\ab[3][1] ), 
	.B(n36), 
	.A(n30));
   NOR2X1M U93 (.Y(\ab[3][0] ), 
	.B(n36), 
	.A(n31));
   NOR2X1M U94 (.Y(\ab[2][7] ), 
	.B(n37), 
	.A(n147));
   NOR2X1M U95 (.Y(\ab[2][6] ), 
	.B(n37), 
	.A(n148));
   NOR2X1M U96 (.Y(\ab[2][5] ), 
	.B(n37), 
	.A(n26));
   NOR2X1M U97 (.Y(\ab[2][4] ), 
	.B(n37), 
	.A(n27));
   NOR2X1M U98 (.Y(\ab[2][3] ), 
	.B(n37), 
	.A(n151));
   NOR2X1M U99 (.Y(\ab[2][2] ), 
	.B(n37), 
	.A(n29));
   NOR2X1M U100 (.Y(\ab[2][1] ), 
	.B(n37), 
	.A(n30));
   NOR2X1M U101 (.Y(\ab[2][0] ), 
	.B(n37), 
	.A(n31));
   NOR2X1M U102 (.Y(\ab[1][7] ), 
	.B(n38), 
	.A(n147));
   NOR2X1M U103 (.Y(\ab[1][6] ), 
	.B(n38), 
	.A(n148));
   NOR2X1M U104 (.Y(\ab[1][5] ), 
	.B(n38), 
	.A(n26));
   NOR2X1M U105 (.Y(\ab[1][4] ), 
	.B(n38), 
	.A(n27));
   NOR2X1M U106 (.Y(\ab[1][3] ), 
	.B(n38), 
	.A(n151));
   NOR2X1M U107 (.Y(\ab[1][2] ), 
	.B(n38), 
	.A(n29));
   NOR2X1M U108 (.Y(\ab[1][1] ), 
	.B(n38), 
	.A(n30));
   NOR2X1M U109 (.Y(\ab[1][0] ), 
	.B(n38), 
	.A(n31));
   NOR2X1M U110 (.Y(\ab[0][7] ), 
	.B(n160), 
	.A(n147));
   NOR2X1M U111 (.Y(\ab[0][6] ), 
	.B(n160), 
	.A(n148));
   NOR2X1M U112 (.Y(\ab[0][5] ), 
	.B(n160), 
	.A(n26));
   NOR2X1M U113 (.Y(\ab[0][4] ), 
	.B(n160), 
	.A(n27));
   NOR2X1M U114 (.Y(\ab[0][3] ), 
	.B(n160), 
	.A(n151));
   NOR2X1M U115 (.Y(\ab[0][2] ), 
	.B(n160), 
	.A(n29));
   NOR2X1M U116 (.Y(\ab[0][1] ), 
	.B(n160), 
	.A(n30));
   NOR2X1M U117 (.Y(PRODUCT[0]), 
	.B(n160), 
	.A(n31));
   ALU_IN_Width8_DW01_add_1 FS_1 (.A({ 1'b0,
		\A1[12] ,
		\A1[11] ,
		\A1[10] ,
		\A1[9] ,
		\A1[8] ,
		\A1[7] ,
		\A1[6] ,
		\SUMB[7][0] ,
		\A1[4] ,
		\A1[3] ,
		\A1[2] ,
		\A1[1] ,
		\A1[0]  }), 
	.B({ n10,
		n14,
		n16,
		n13,
		n15,
		n12,
		n11,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }), 
	.CI(1'b0), 
	.SUM({ PRODUCT[15],
		PRODUCT[14],
		PRODUCT[13],
		PRODUCT[12],
		PRODUCT[11],
		PRODUCT[10],
		PRODUCT[9],
		PRODUCT[8],
		PRODUCT[7],
		PRODUCT[6],
		PRODUCT[5],
		PRODUCT[4],
		PRODUCT[3],
		PRODUCT[2] }));
endmodule

module ALU_IN_Width8_test_1 (
	CLK, 
	RST, 
	EN, 
	ALU_FUN, 
	A, 
	B, 
	ALU_OUT, 
	OUT_Valid, 
	test_si2, 
	test_si1, 
	test_se, 
	FE_OFN4_M_Domain1_SYNC_RST);
   input CLK;
   input RST;
   input EN;
   input [3:0] ALU_FUN;
   input [7:0] A;
   input [7:0] B;
   output [15:0] ALU_OUT;
   output OUT_Valid;
   input test_si2;
   input test_si1;
   input test_se;
   input FE_OFN4_M_Domain1_SYNC_RST;

   // Internal wires
   wire FE_OFN6_n57;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N124;
   wire N125;
   wire N127;
   wire N128;
   wire N129;
   wire N130;
   wire N131;
   wire N132;
   wire N133;
   wire N134;
   wire N167;
   wire N168;
   wire N169;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n3;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire [15:0] Com_ALU_OUT;

   BUFX2M FE_OFC6_n57 (.Y(FE_OFN6_n57), 
	.A(n57));
   SDFFRQX2M \ALU_OUT_reg[15]  (.SI(ALU_OUT[14]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(ALU_OUT[15]), 
	.D(Com_ALU_OUT[15]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[14]  (.SI(ALU_OUT[13]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(ALU_OUT[14]), 
	.D(Com_ALU_OUT[14]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[13]  (.SI(ALU_OUT[12]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(ALU_OUT[13]), 
	.D(Com_ALU_OUT[13]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[12]  (.SI(ALU_OUT[11]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(ALU_OUT[12]), 
	.D(Com_ALU_OUT[12]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[11]  (.SI(ALU_OUT[10]), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(ALU_OUT[11]), 
	.D(Com_ALU_OUT[11]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[10]  (.SI(ALU_OUT[9]), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(ALU_OUT[10]), 
	.D(Com_ALU_OUT[10]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[9]  (.SI(ALU_OUT[8]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(ALU_OUT[9]), 
	.D(Com_ALU_OUT[9]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[8]  (.SI(test_si2), 
	.SE(test_se), 
	.RN(RST), 
	.Q(ALU_OUT[8]), 
	.D(Com_ALU_OUT[8]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[7]  (.SI(ALU_OUT[6]), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(ALU_OUT[7]), 
	.D(Com_ALU_OUT[7]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[6]  (.SI(ALU_OUT[5]), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(ALU_OUT[6]), 
	.D(Com_ALU_OUT[6]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[5]  (.SI(ALU_OUT[4]), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(ALU_OUT[5]), 
	.D(Com_ALU_OUT[5]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[4]  (.SI(ALU_OUT[3]), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(ALU_OUT[4]), 
	.D(Com_ALU_OUT[4]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[3]  (.SI(ALU_OUT[2]), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(ALU_OUT[3]), 
	.D(Com_ALU_OUT[3]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[2]  (.SI(ALU_OUT[1]), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(ALU_OUT[2]), 
	.D(Com_ALU_OUT[2]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[1]  (.SI(ALU_OUT[0]), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(ALU_OUT[1]), 
	.D(Com_ALU_OUT[1]), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[0]  (.SI(test_si1), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(ALU_OUT[0]), 
	.D(Com_ALU_OUT[0]), 
	.CK(CLK));
   SDFFRQX2M OUT_Valid_reg (.SI(ALU_OUT[15]), 
	.SE(test_se), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(OUT_Valid), 
	.D(EN), 
	.CK(CLK));
   INVX2M U26 (.Y(n164), 
	.A(n70));
   INVX2M U27 (.Y(n163), 
	.A(n114));
   INVX2M U28 (.Y(n162), 
	.A(n64));
   INVX2M U29 (.Y(n161), 
	.A(n119));
   OAI2BB1X2M U30 (.Y(Com_ALU_OUT[9]), 
	.B0(n53), 
	.A1N(n52), 
	.A0N(N119));
   OAI2BB1X2M U31 (.Y(Com_ALU_OUT[10]), 
	.B0(n53), 
	.A1N(n52), 
	.A0N(N120));
   OAI2BB1X2M U32 (.Y(Com_ALU_OUT[11]), 
	.B0(n53), 
	.A1N(n52), 
	.A0N(N121));
   OAI2BB1X2M U33 (.Y(Com_ALU_OUT[12]), 
	.B0(n53), 
	.A1N(n52), 
	.A0N(N122));
   OAI2BB1X2M U34 (.Y(Com_ALU_OUT[13]), 
	.B0(n53), 
	.A1N(n52), 
	.A0N(N123));
   OAI2BB1X2M U35 (.Y(Com_ALU_OUT[14]), 
	.B0(n53), 
	.A1N(n52), 
	.A0N(N124));
   OAI2BB1X2M U36 (.Y(Com_ALU_OUT[15]), 
	.B0(n53), 
	.A1N(n52), 
	.A0N(N125));
   OAI2B11X2M U37 (.Y(n59), 
	.C0(n163), 
	.B0(n164), 
	.A1N(N109), 
	.A0(n119));
   OAI21X2M U38 (.Y(n69), 
	.B0(n128), 
	.A1(n129), 
	.A0(n3));
   NOR2X2M U39 (.Y(n70), 
	.B(n3), 
	.A(n118));
   NOR2BX2M U40 (.Y(n58), 
	.B(n3), 
	.AN(n130));
   OAI2B1X2M U41 (.Y(n114), 
	.B0(n128), 
	.A1N(n127), 
	.A0(n118));
   NAND2X2M U42 (.Y(n53), 
	.B(n59), 
	.A(EN));
   OAI2BB2X1M U43 (.Y(n63), 
	.B1(n64), 
	.B0(n154), 
	.A1N(FE_OFN6_n57), 
	.A0N(N117));
   NAND2X2M U44 (.Y(n64), 
	.B(n127), 
	.A(n166));
   NOR2BX2M U45 (.Y(n52), 
	.B(n169), 
	.AN(FE_OFN6_n57));
   NAND2X2M U46 (.Y(n119), 
	.B(n127), 
	.A(n130));
   INVX2M U47 (.Y(n165), 
	.A(n67));
   INVX2M U48 (.Y(n166), 
	.A(n129));
   INVX2M U49 (.Y(n169), 
	.A(EN));
   NOR3BX2M U50 (.Y(n56), 
	.C(ALU_FUN[0]), 
	.B(n118), 
	.AN(ALU_FUN[3]));
   NOR3BX2M U51 (.Y(n74), 
	.C(n129), 
	.B(n168), 
	.AN(ALU_FUN[3]));
   NOR3X2M U52 (.Y(n57), 
	.C(n167), 
	.B(ALU_FUN[2]), 
	.A(n3));
   OAI221X1M U53 (.Y(n106), 
	.C0(n164), 
	.B1(n159), 
	.B0(n67), 
	.A1(n163), 
	.A0(A[2]));
   OAI221X1M U54 (.Y(n99), 
	.C0(n164), 
	.B1(n158), 
	.B0(n67), 
	.A1(n163), 
	.A0(A[3]));
   OAI221X1M U55 (.Y(n92), 
	.C0(n164), 
	.B1(n157), 
	.B0(n67), 
	.A1(n163), 
	.A0(A[4]));
   OAI221X1M U56 (.Y(n85), 
	.C0(n164), 
	.B1(n156), 
	.B0(n67), 
	.A1(n163), 
	.A0(A[5]));
   OAI221X1M U57 (.Y(n78), 
	.C0(n164), 
	.B1(n155), 
	.B0(n67), 
	.A1(n163), 
	.A0(A[6]));
   OAI221X1M U58 (.Y(n66), 
	.C0(n164), 
	.B1(n67), 
	.B0(n154), 
	.A1(n163), 
	.A0(A[7]));
   NOR2X2M U59 (.Y(n130), 
	.B(ALU_FUN[1]), 
	.A(ALU_FUN[2]));
   INVX2M U60 (.Y(n145), 
	.A(n33));
   NOR2X2M U61 (.Y(n127), 
	.B(ALU_FUN[3]), 
	.A(n168));
   OAI2B2X1M U62 (.Y(n111), 
	.B1(n113), 
	.B0(B[1]), 
	.A1N(B[1]), 
	.A0(n112));
   AOI221XLM U63 (.Y(n112), 
	.C0(n162), 
	.B1(n69), 
	.B0(A[1]), 
	.A1(n143), 
	.A0(n165));
   AOI221XLM U64 (.Y(n113), 
	.C0(n70), 
	.B1(n143), 
	.B0(n114), 
	.A1(n165), 
	.A0(A[1]));
   NAND2X2M U65 (.Y(n118), 
	.B(ALU_FUN[1]), 
	.A(ALU_FUN[2]));
   NAND2X2M U66 (.Y(n129), 
	.B(n167), 
	.A(ALU_FUN[2]));
   NOR3X2M U67 (.Y(n132), 
	.C(ALU_FUN[0]), 
	.B(ALU_FUN[2]), 
	.A(n167));
   INVX2M U68 (.Y(n168), 
	.A(ALU_FUN[0]));
   INVX2M U69 (.Y(n167), 
	.A(ALU_FUN[1]));
   NAND3X2M U70 (.Y(n67), 
	.C(ALU_FUN[3]), 
	.B(n168), 
	.A(n130));
   NAND3X2M U71 (.Y(n128), 
	.C(ALU_FUN[3]), 
	.B(ALU_FUN[0]), 
	.A(n130));
   AOI31X2M U72 (.Y(Com_ALU_OUT[4]), 
	.B0(n169), 
	.A2(n88), 
	.A1(n87), 
	.A0(n86));
   AOI22X1M U73 (.Y(n86), 
	.B1(n58), 
	.B0(N96), 
	.A1(n161), 
	.A0(N105));
   AOI221XLM U74 (.Y(n88), 
	.C0(n89), 
	.B1(A[5]), 
	.B0(n74), 
	.A1(n56), 
	.A0(A[3]));
   AOI222X1M U75 (.Y(n87), 
	.C1(n162), 
	.C0(A[4]), 
	.B1(n157), 
	.B0(n70), 
	.A1(FE_OFN6_n57), 
	.A0(N114));
   AOI31X2M U76 (.Y(Com_ALU_OUT[5]), 
	.B0(n169), 
	.A2(n81), 
	.A1(n80), 
	.A0(n79));
   AOI22X1M U77 (.Y(n79), 
	.B1(n58), 
	.B0(N97), 
	.A1(n161), 
	.A0(N106));
   AOI221XLM U78 (.Y(n81), 
	.C0(n82), 
	.B1(A[6]), 
	.B0(n74), 
	.A1(n56), 
	.A0(A[4]));
   AOI222X1M U79 (.Y(n80), 
	.C1(n162), 
	.C0(A[5]), 
	.B1(n156), 
	.B0(n70), 
	.A1(FE_OFN6_n57), 
	.A0(N115));
   AOI31X2M U80 (.Y(Com_ALU_OUT[6]), 
	.B0(n169), 
	.A2(n73), 
	.A1(n72), 
	.A0(n71));
   AOI22X1M U81 (.Y(n71), 
	.B1(n58), 
	.B0(N98), 
	.A1(n161), 
	.A0(N107));
   AOI221XLM U82 (.Y(n73), 
	.C0(n75), 
	.B1(A[7]), 
	.B0(n74), 
	.A1(n56), 
	.A0(A[5]));
   AOI222X1M U83 (.Y(n72), 
	.C1(A[6]), 
	.C0(n162), 
	.B1(n155), 
	.B0(n70), 
	.A1(FE_OFN6_n57), 
	.A0(N116));
   AOI31X2M U84 (.Y(Com_ALU_OUT[2]), 
	.B0(n169), 
	.A2(n102), 
	.A1(n101), 
	.A0(n100));
   AOI22X1M U85 (.Y(n100), 
	.B1(n58), 
	.B0(N94), 
	.A1(n161), 
	.A0(N103));
   AOI221XLM U86 (.Y(n102), 
	.C0(n103), 
	.B1(n74), 
	.B0(A[3]), 
	.A1(n56), 
	.A0(A[1]));
   AOI222X1M U87 (.Y(n101), 
	.C1(n162), 
	.C0(A[2]), 
	.B1(n159), 
	.B0(n70), 
	.A1(FE_OFN6_n57), 
	.A0(N112));
   AOI31X2M U88 (.Y(Com_ALU_OUT[3]), 
	.B0(n169), 
	.A2(n95), 
	.A1(n94), 
	.A0(n93));
   AOI22X1M U89 (.Y(n93), 
	.B1(n58), 
	.B0(N95), 
	.A1(n161), 
	.A0(N104));
   AOI221XLM U90 (.Y(n95), 
	.C0(n96), 
	.B1(n74), 
	.B0(A[4]), 
	.A1(n56), 
	.A0(A[2]));
   AOI222X1M U91 (.Y(n94), 
	.C1(n162), 
	.C0(A[3]), 
	.B1(n158), 
	.B0(n70), 
	.A1(FE_OFN6_n57), 
	.A0(N113));
   AOI31X2M U92 (.Y(Com_ALU_OUT[0]), 
	.B0(n169), 
	.A2(n122), 
	.A1(n121), 
	.A0(n120));
   AOI22X1M U93 (.Y(n120), 
	.B1(n58), 
	.B0(N92), 
	.A1(n161), 
	.A0(N101));
   AOI211X2M U94 (.Y(n122), 
	.C0(n124), 
	.B0(n123), 
	.A1(n74), 
	.A0(A[1]));
   AOI222X1M U95 (.Y(n121), 
	.C1(n162), 
	.C0(A[0]), 
	.B1(n160), 
	.B0(n70), 
	.A1(FE_OFN6_n57), 
	.A0(N110));
   AOI31X2M U96 (.Y(Com_ALU_OUT[1]), 
	.B0(n169), 
	.A2(n109), 
	.A1(n108), 
	.A0(n107));
   AOI211X2M U97 (.Y(n109), 
	.C0(n111), 
	.B0(n110), 
	.A1(n56), 
	.A0(A[0]));
   AOI222X1M U98 (.Y(n108), 
	.C1(n143), 
	.C0(n70), 
	.B1(n74), 
	.B0(A[2]), 
	.A1(n162), 
	.A0(A[1]));
   AOI222X1M U99 (.Y(n107), 
	.C1(n161), 
	.C0(N102), 
	.B1(FE_OFN6_n57), 
	.B0(N111), 
	.A1(n58), 
	.A0(N93));
   AOI31X2M U100 (.Y(Com_ALU_OUT[7]), 
	.B0(n169), 
	.A2(n62), 
	.A1(n61), 
	.A0(n60));
   AOI22X1M U101 (.Y(n60), 
	.B1(n154), 
	.B0(n70), 
	.A1(n56), 
	.A0(A[6]));
   AOI221XLM U102 (.Y(n62), 
	.C0(n63), 
	.B1(n58), 
	.B0(N99), 
	.A1(n161), 
	.A0(N108));
   AOI222X1M U103 (.Y(n61), 
	.C1(n147), 
	.C0(n66), 
	.B1(n65), 
	.B0(N134), 
	.A1(n153), 
	.A0(B[7]));
   INVX2M U104 (.Y(n146), 
	.A(n44));
   OAI21X2M U105 (.Y(n75), 
	.B0(n77), 
	.A1(n148), 
	.A0(n76));
   AOI22X1M U106 (.Y(n77), 
	.B1(n148), 
	.B0(n78), 
	.A1(n65), 
	.A0(N133));
   AOI221XLM U107 (.Y(n76), 
	.C0(n162), 
	.B1(n69), 
	.B0(A[6]), 
	.A1(n155), 
	.A0(n165));
   INVX2M U108 (.Y(n148), 
	.A(B[6]));
   AOI21X2M U109 (.Y(Com_ALU_OUT[8]), 
	.B0(n169), 
	.A1(n55), 
	.A0(n54));
   AOI21X2M U110 (.Y(n54), 
	.B0(n59), 
	.A1(n58), 
	.A0(N100));
   AOI22X1M U111 (.Y(n55), 
	.B1(FE_OFN6_n57), 
	.B0(N118), 
	.A1(n56), 
	.A0(A[7]));
   OR2X2M U112 (.Y(n3), 
	.B(ALU_FUN[0]), 
	.A(ALU_FUN[3]));
   INVX2M U113 (.Y(n153), 
	.A(n68));
   AOI221XLM U114 (.Y(n68), 
	.C0(n162), 
	.B1(n165), 
	.B0(n154), 
	.A1(A[7]), 
	.A0(n69));
   OAI2BB1X2M U115 (.Y(n123), 
	.B0(n131), 
	.A1N(n65), 
	.A0N(N127));
   AOI31X2M U116 (.Y(n131), 
	.B0(n117), 
	.A2(n132), 
	.A1(ALU_FUN[3]), 
	.A0(N167));
   AND4X2M U117 (.Y(n117), 
	.D(n168), 
	.C(ALU_FUN[3]), 
	.B(n166), 
	.A(N169));
   OAI2BB1X2M U118 (.Y(n110), 
	.B0(n115), 
	.A1N(n65), 
	.A0N(N128));
   AOI31X2M U119 (.Y(n115), 
	.B0(n117), 
	.A2(n116), 
	.A1(ALU_FUN[3]), 
	.A0(N168));
   NOR3X2M U120 (.Y(n116), 
	.C(n167), 
	.B(ALU_FUN[2]), 
	.A(n168));
   INVX2M U121 (.Y(n154), 
	.A(A[7]));
   INVX2M U122 (.Y(n155), 
	.A(A[6]));
   INVX2M U123 (.Y(n160), 
	.A(A[0]));
   INVX2M U124 (.Y(n159), 
	.A(A[2]));
   INVX2M U125 (.Y(n158), 
	.A(A[3]));
   INVX2M U126 (.Y(n156), 
	.A(A[5]));
   INVX2M U127 (.Y(n157), 
	.A(A[4]));
   INVX2M U128 (.Y(n143), 
	.A(A[1]));
   INVX2M U129 (.Y(n147), 
	.A(B[7]));
   OAI2B2X1M U130 (.Y(n124), 
	.B1(n126), 
	.B0(B[0]), 
	.A1N(B[0]), 
	.A0(n125));
   AOI221XLM U131 (.Y(n125), 
	.C0(n162), 
	.B1(n69), 
	.B0(A[0]), 
	.A1(n160), 
	.A0(n165));
   AOI221XLM U132 (.Y(n126), 
	.C0(n70), 
	.B1(n160), 
	.B0(n114), 
	.A1(n165), 
	.A0(A[0]));
   AND3X2M U133 (.Y(n65), 
	.C(n133), 
	.B(ALU_FUN[1]), 
	.A(n127));
   AOI21X2M U134 (.Y(n133), 
	.B0(ALU_FUN[2]), 
	.A1(n135), 
	.A0(n134));
   NOR4X1M U135 (.Y(n135), 
	.D(B[4]), 
	.C(B[5]), 
	.B(B[6]), 
	.A(B[7]));
   NOR4X1M U136 (.Y(n134), 
	.D(B[0]), 
	.C(B[1]), 
	.B(B[2]), 
	.A(B[3]));
   OAI21X2M U137 (.Y(n103), 
	.B0(n105), 
	.A1(n152), 
	.A0(n104));
   AOI22X1M U138 (.Y(n105), 
	.B1(n152), 
	.B0(n106), 
	.A1(n65), 
	.A0(N129));
   AOI221XLM U139 (.Y(n104), 
	.C0(n162), 
	.B1(n69), 
	.B0(A[2]), 
	.A1(n159), 
	.A0(n165));
   INVX2M U140 (.Y(n152), 
	.A(B[2]));
   OAI21X2M U141 (.Y(n96), 
	.B0(n98), 
	.A1(n151), 
	.A0(n97));
   AOI22X1M U142 (.Y(n98), 
	.B1(n151), 
	.B0(n99), 
	.A1(n65), 
	.A0(N130));
   AOI221XLM U143 (.Y(n97), 
	.C0(n162), 
	.B1(n69), 
	.B0(A[3]), 
	.A1(n158), 
	.A0(n165));
   INVX2M U144 (.Y(n151), 
	.A(B[3]));
   OAI21X2M U145 (.Y(n89), 
	.B0(n91), 
	.A1(n150), 
	.A0(n90));
   AOI22X1M U146 (.Y(n91), 
	.B1(n150), 
	.B0(n92), 
	.A1(n65), 
	.A0(N131));
   AOI221XLM U147 (.Y(n90), 
	.C0(n162), 
	.B1(n69), 
	.B0(A[4]), 
	.A1(n157), 
	.A0(n165));
   INVX2M U148 (.Y(n150), 
	.A(B[4]));
   OAI21X2M U149 (.Y(n82), 
	.B0(n84), 
	.A1(n149), 
	.A0(n83));
   AOI22X1M U150 (.Y(n84), 
	.B1(n149), 
	.B0(n85), 
	.A1(n65), 
	.A0(N132));
   AOI221XLM U151 (.Y(n83), 
	.C0(n162), 
	.B1(n69), 
	.B0(A[5]), 
	.A1(n156), 
	.A0(n165));
   INVX2M U152 (.Y(n149), 
	.A(B[5]));
   INVX2M U161 (.Y(n144), 
	.A(B[0]));
   NOR2X1M U162 (.Y(n139), 
	.B(B[7]), 
	.A(n154));
   NAND2BX1M U163 (.Y(n48), 
	.B(A[4]), 
	.AN(B[4]));
   NAND2BX1M U164 (.Y(n37), 
	.B(B[4]), 
	.AN(A[4]));
   CLKNAND2X2M U165 (.Y(n50), 
	.B(n37), 
	.A(n48));
   NOR2X1M U166 (.Y(n45), 
	.B(A[3]), 
	.A(n151));
   NOR2X1M U167 (.Y(n36), 
	.B(A[2]), 
	.A(n152));
   NOR2X1M U168 (.Y(n33), 
	.B(A[0]), 
	.A(n144));
   CLKNAND2X2M U169 (.Y(n47), 
	.B(n152), 
	.A(A[2]));
   NAND2BX1M U170 (.Y(n42), 
	.B(n47), 
	.AN(n36));
   AOI21X1M U171 (.Y(n34), 
	.B0(B[1]), 
	.A1(n143), 
	.A0(n33));
   AOI211X1M U172 (.Y(n35), 
	.C0(n34), 
	.B0(n42), 
	.A1(n145), 
	.A0(A[1]));
   CLKNAND2X2M U173 (.Y(n46), 
	.B(n151), 
	.A(A[3]));
   OAI31X1M U174 (.Y(n38), 
	.B0(n46), 
	.A2(n35), 
	.A1(n36), 
	.A0(n45));
   NAND2BX1M U175 (.Y(n137), 
	.B(B[5]), 
	.AN(A[5]));
   OAI211X1M U176 (.Y(n39), 
	.C0(n137), 
	.B0(n37), 
	.A1(n38), 
	.A0(n50));
   NAND2BX1M U177 (.Y(n49), 
	.B(A[5]), 
	.AN(B[5]));
   XNOR2X1M U178 (.Y(n136), 
	.B(B[6]), 
	.A(A[6]));
   AOI32X1M U179 (.Y(n40), 
	.B1(n155), 
	.B0(B[6]), 
	.A2(n136), 
	.A1(n49), 
	.A0(n39));
   CLKNAND2X2M U180 (.Y(n140), 
	.B(n154), 
	.A(B[7]));
   OAI21X1M U181 (.Y(N169), 
	.B0(n140), 
	.A1(n40), 
	.A0(n139));
   CLKNAND2X2M U182 (.Y(n43), 
	.B(n144), 
	.A(A[0]));
   OA21X1M U183 (.Y(n41), 
	.B0(B[1]), 
	.A1(n143), 
	.A0(n43));
   AOI211X1M U184 (.Y(n44), 
	.C0(n41), 
	.B0(n42), 
	.A1(n143), 
	.A0(n43));
   AOI31X1M U185 (.Y(n51), 
	.B0(n45), 
	.A2(n46), 
	.A1(n47), 
	.A0(n146));
   OAI2B11X1M U186 (.Y(n138), 
	.C0(n48), 
	.B0(n49), 
	.A1N(n51), 
	.A0(n50));
   AOI32X1M U187 (.Y(n141), 
	.B1(n148), 
	.B0(A[6]), 
	.A2(n136), 
	.A1(n137), 
	.A0(n138));
   AOI2B1X1M U188 (.Y(n142), 
	.B0(n139), 
	.A1N(n141), 
	.A0(n140));
   CLKINVX1M U189 (.Y(N168), 
	.A(n142));
   NOR2X1M U190 (.Y(N167), 
	.B(N168), 
	.A(N169));
   ALU_IN_Width8_DW_div_uns_0 div_51 (.a({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }), 
	.b({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }), 
	.quotient({ N134,
		N133,
		N132,
		N131,
		N130,
		N129,
		N128,
		N127 }), 
	.n144(n144), 
	.n151(n151), 
	.n152(n152), 
	.n149(n149), 
	.n150(n150), 
	.n160(n160), 
	.n143(n143), 
	.n159(n159), 
	.n158(n158), 
	.n157(n157), 
	.n156(n156), 
	.n155(n155), 
	.n148(n148), 
	.n147(n147));
   ALU_IN_Width8_DW01_sub_0 sub_43 (.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }), 
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }), 
	.CI(1'b0), 
	.DIFF({ N109,
		N108,
		N107,
		N106,
		N105,
		N104,
		N103,
		N102,
		N101 }), 
	.n144(n144), 
	.n151(n151), 
	.n152(n152), 
	.n149(n149), 
	.n150(n150), 
	.n160(n160), 
	.n148(n148), 
	.n147(n147));
   ALU_IN_Width8_DW01_add_0 add_39 (.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }), 
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }), 
	.CI(1'b0), 
	.SUM({ N100,
		N99,
		N98,
		N97,
		N96,
		N95,
		N94,
		N93,
		N92 }));
   ALU_IN_Width8_DW02_mult_0 mult_47 (.A({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }), 
	.B({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }), 
	.TC(1'b0), 
	.PRODUCT({ N125,
		N124,
		N123,
		N122,
		N121,
		N120,
		N119,
		N118,
		N117,
		N116,
		N115,
		N114,
		N113,
		N112,
		N111,
		N110 }), 
	.n144(n144), 
	.n151(n151), 
	.n152(n152), 
	.n149(n149), 
	.n150(n150), 
	.n160(n160), 
	.n143(n143), 
	.n159(n159), 
	.n158(n158), 
	.n157(n157), 
	.n156(n156), 
	.n155(n155), 
	.n154(n154), 
	.n148(n148), 
	.n147(n147));
endmodule

module Reg_File_WIDTH8_DEPTH16_ADDR4_test_1 (
	CLK, 
	RST, 
	WrEn, 
	RdEn, 
	Address, 
	WrData, 
	RdData, 
	RdData_VLD, 
	REG0, 
	REG1, 
	REG2, 
	REG3, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN2_M_Domain1_SYNC_RST, 
	FE_OFN4_M_Domain1_SYNC_RST, 
	REF_CLK_M__L5_N11, 
	REF_CLK_M__L5_N12, 
	REF_CLK_M__L5_N13, 
	REF_CLK_M__L5_N14, 
	REF_CLK_M__L5_N15, 
	REF_CLK_M__L5_N3, 
	REF_CLK_M__L5_N8, 
	REF_CLK_M__L5_N9);
   input CLK;
   input RST;
   input WrEn;
   input RdEn;
   input [3:0] Address;
   input [7:0] WrData;
   output [7:0] RdData;
   output RdData_VLD;
   output [7:0] REG0;
   output [7:0] REG1;
   output [7:0] REG2;
   output [7:0] REG3;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN2_M_Domain1_SYNC_RST;
   input FE_OFN4_M_Domain1_SYNC_RST;
   input REF_CLK_M__L5_N11;
   input REF_CLK_M__L5_N12;
   input REF_CLK_M__L5_N13;
   input REF_CLK_M__L5_N14;
   input REF_CLK_M__L5_N15;
   input REF_CLK_M__L5_N3;
   input REF_CLK_M__L5_N8;
   input REF_CLK_M__L5_N9;

   // Internal wires
   wire FE_OFN3_M_Domain1_SYNC_RST;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire \memory[15][7] ;
   wire \memory[15][6] ;
   wire \memory[15][5] ;
   wire \memory[15][4] ;
   wire \memory[15][3] ;
   wire \memory[15][2] ;
   wire \memory[15][1] ;
   wire \memory[15][0] ;
   wire \memory[14][7] ;
   wire \memory[14][6] ;
   wire \memory[14][5] ;
   wire \memory[14][4] ;
   wire \memory[14][3] ;
   wire \memory[14][2] ;
   wire \memory[14][1] ;
   wire \memory[14][0] ;
   wire \memory[13][7] ;
   wire \memory[13][6] ;
   wire \memory[13][5] ;
   wire \memory[13][4] ;
   wire \memory[13][3] ;
   wire \memory[13][2] ;
   wire \memory[13][1] ;
   wire \memory[13][0] ;
   wire \memory[12][7] ;
   wire \memory[12][6] ;
   wire \memory[12][5] ;
   wire \memory[12][4] ;
   wire \memory[12][3] ;
   wire \memory[12][2] ;
   wire \memory[12][1] ;
   wire \memory[12][0] ;
   wire \memory[11][7] ;
   wire \memory[11][6] ;
   wire \memory[11][5] ;
   wire \memory[11][4] ;
   wire \memory[11][3] ;
   wire \memory[11][2] ;
   wire \memory[11][1] ;
   wire \memory[11][0] ;
   wire \memory[10][7] ;
   wire \memory[10][6] ;
   wire \memory[10][5] ;
   wire \memory[10][4] ;
   wire \memory[10][3] ;
   wire \memory[10][2] ;
   wire \memory[10][1] ;
   wire \memory[10][0] ;
   wire \memory[9][7] ;
   wire \memory[9][6] ;
   wire \memory[9][5] ;
   wire \memory[9][4] ;
   wire \memory[9][3] ;
   wire \memory[9][2] ;
   wire \memory[9][1] ;
   wire \memory[9][0] ;
   wire \memory[8][7] ;
   wire \memory[8][6] ;
   wire \memory[8][5] ;
   wire \memory[8][4] ;
   wire \memory[8][3] ;
   wire \memory[8][2] ;
   wire \memory[8][1] ;
   wire \memory[8][0] ;
   wire \memory[7][7] ;
   wire \memory[7][6] ;
   wire \memory[7][5] ;
   wire \memory[7][4] ;
   wire \memory[7][3] ;
   wire \memory[7][2] ;
   wire \memory[7][1] ;
   wire \memory[7][0] ;
   wire \memory[6][7] ;
   wire \memory[6][6] ;
   wire \memory[6][5] ;
   wire \memory[6][4] ;
   wire \memory[6][3] ;
   wire \memory[6][2] ;
   wire \memory[6][1] ;
   wire \memory[6][0] ;
   wire \memory[5][7] ;
   wire \memory[5][6] ;
   wire \memory[5][5] ;
   wire \memory[5][4] ;
   wire \memory[5][3] ;
   wire \memory[5][2] ;
   wire \memory[5][1] ;
   wire \memory[5][0] ;
   wire \memory[4][7] ;
   wire \memory[4][6] ;
   wire \memory[4][5] ;
   wire \memory[4][4] ;
   wire \memory[4][3] ;
   wire \memory[4][2] ;
   wire \memory[4][1] ;
   wire \memory[4][0] ;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n336;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n370;
   wire n371;
   wire n372;
   wire n373;

   assign N11 = Address[0] ;
   assign N12 = Address[1] ;
   assign N13 = Address[2] ;
   assign N14 = Address[3] ;
   assign test_so2 = \memory[15][7]  ;
   assign test_so1 = \memory[8][6]  ;

   CLKINVX6M FE_OFC3_M_Domain1_SYNC_RST (.Y(FE_OFN3_M_Domain1_SYNC_RST), 
	.A(RST));
   SDFFRQX2M \memory_reg[13][7]  (.SI(\memory[13][6] ), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[13][7] ), 
	.D(n298), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[13][6]  (.SI(\memory[13][5] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[13][6] ), 
	.D(n297), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[13][5]  (.SI(\memory[13][4] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[13][5] ), 
	.D(n296), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[13][4]  (.SI(\memory[13][3] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[13][4] ), 
	.D(n295), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[13][3]  (.SI(\memory[13][2] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[13][3] ), 
	.D(n294), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[13][2]  (.SI(\memory[13][1] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[13][2] ), 
	.D(n293), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[13][1]  (.SI(\memory[13][0] ), 
	.SE(n371), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[13][1] ), 
	.D(n292), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[13][0]  (.SI(\memory[12][7] ), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[13][0] ), 
	.D(n291), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[9][7]  (.SI(\memory[9][6] ), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[9][7] ), 
	.D(n266), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[9][6]  (.SI(\memory[9][5] ), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[9][6] ), 
	.D(n265), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[9][5]  (.SI(\memory[9][4] ), 
	.SE(n371), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[9][5] ), 
	.D(n264), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[9][4]  (.SI(\memory[9][3] ), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[9][4] ), 
	.D(n263), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[9][3]  (.SI(\memory[9][2] ), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[9][3] ), 
	.D(n262), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[9][2]  (.SI(\memory[9][1] ), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[9][2] ), 
	.D(n261), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[9][1]  (.SI(\memory[9][0] ), 
	.SE(n371), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[9][1] ), 
	.D(n260), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[9][0]  (.SI(\memory[8][7] ), 
	.SE(n370), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(\memory[9][0] ), 
	.D(n259), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[5][7]  (.SI(\memory[5][6] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[5][7] ), 
	.D(n234), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[5][6]  (.SI(\memory[5][5] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[5][6] ), 
	.D(n233), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[5][5]  (.SI(\memory[5][4] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[5][5] ), 
	.D(n232), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[5][4]  (.SI(\memory[5][3] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[5][4] ), 
	.D(n231), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[5][3]  (.SI(\memory[5][2] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[5][3] ), 
	.D(n230), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[5][2]  (.SI(\memory[5][1] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[5][2] ), 
	.D(n229), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[5][1]  (.SI(\memory[5][0] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[5][1] ), 
	.D(n228), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[5][0]  (.SI(\memory[4][7] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[5][0] ), 
	.D(n227), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[15][7]  (.SI(\memory[15][6] ), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[15][7] ), 
	.D(n314), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[15][6]  (.SI(\memory[15][5] ), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[15][6] ), 
	.D(n313), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[15][5]  (.SI(\memory[15][4] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[15][5] ), 
	.D(n312), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[15][4]  (.SI(\memory[15][3] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[15][4] ), 
	.D(n311), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[15][3]  (.SI(\memory[15][2] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[15][3] ), 
	.D(n310), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[15][2]  (.SI(\memory[15][1] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[15][2] ), 
	.D(n309), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[15][1]  (.SI(\memory[15][0] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[15][1] ), 
	.D(n308), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[15][0]  (.SI(\memory[14][7] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[15][0] ), 
	.D(n307), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[11][7]  (.SI(\memory[11][6] ), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[11][7] ), 
	.D(n282), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[11][6]  (.SI(\memory[11][5] ), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[11][6] ), 
	.D(n281), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[11][5]  (.SI(\memory[11][4] ), 
	.SE(n371), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[11][5] ), 
	.D(n280), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[11][4]  (.SI(\memory[11][3] ), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[11][4] ), 
	.D(n279), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[11][3]  (.SI(\memory[11][2] ), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[11][3] ), 
	.D(n278), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[11][2]  (.SI(\memory[11][1] ), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[11][2] ), 
	.D(n277), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[11][1]  (.SI(\memory[11][0] ), 
	.SE(n371), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[11][1] ), 
	.D(n276), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[11][0]  (.SI(\memory[10][7] ), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[11][0] ), 
	.D(n275), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[7][7]  (.SI(\memory[7][6] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[7][7] ), 
	.D(n250), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[7][6]  (.SI(\memory[7][5] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[7][6] ), 
	.D(n249), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[7][5]  (.SI(\memory[7][4] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[7][5] ), 
	.D(n248), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[7][4]  (.SI(\memory[7][3] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[7][4] ), 
	.D(n247), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[7][3]  (.SI(\memory[7][2] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[7][3] ), 
	.D(n246), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[7][2]  (.SI(\memory[7][1] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[7][2] ), 
	.D(n245), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[7][1]  (.SI(\memory[7][0] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[7][1] ), 
	.D(n244), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[7][0]  (.SI(\memory[6][7] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[7][0] ), 
	.D(n243), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \memory_reg[14][7]  (.SI(\memory[14][6] ), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[14][7] ), 
	.D(n306), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[14][6]  (.SI(\memory[14][5] ), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[14][6] ), 
	.D(n305), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[14][5]  (.SI(\memory[14][4] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[14][5] ), 
	.D(n304), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[14][4]  (.SI(\memory[14][3] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[14][4] ), 
	.D(n303), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[14][3]  (.SI(\memory[14][2] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[14][3] ), 
	.D(n302), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[14][2]  (.SI(\memory[14][1] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[14][2] ), 
	.D(n301), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[14][1]  (.SI(\memory[14][0] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[14][1] ), 
	.D(n300), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[14][0]  (.SI(\memory[13][7] ), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[14][0] ), 
	.D(n299), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[10][7]  (.SI(\memory[10][6] ), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[10][7] ), 
	.D(n274), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[10][6]  (.SI(\memory[10][5] ), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[10][6] ), 
	.D(n273), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[10][5]  (.SI(\memory[10][4] ), 
	.SE(n371), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[10][5] ), 
	.D(n272), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[10][4]  (.SI(\memory[10][3] ), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[10][4] ), 
	.D(n271), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[10][3]  (.SI(\memory[10][2] ), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[10][3] ), 
	.D(n270), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[10][2]  (.SI(\memory[10][1] ), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[10][2] ), 
	.D(n269), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[10][1]  (.SI(\memory[10][0] ), 
	.SE(n371), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[10][1] ), 
	.D(n268), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[10][0]  (.SI(\memory[9][7] ), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[10][0] ), 
	.D(n267), 
	.CK(REF_CLK_M__L5_N11));
   SDFFRQX2M \memory_reg[6][7]  (.SI(\memory[6][6] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[6][7] ), 
	.D(n242), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[6][6]  (.SI(\memory[6][5] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[6][6] ), 
	.D(n241), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[6][5]  (.SI(\memory[6][4] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[6][5] ), 
	.D(n240), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[6][4]  (.SI(\memory[6][3] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[6][4] ), 
	.D(n239), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[6][3]  (.SI(\memory[6][2] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[6][3] ), 
	.D(n238), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[6][2]  (.SI(\memory[6][1] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[6][2] ), 
	.D(n237), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \memory_reg[6][1]  (.SI(\memory[6][0] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[6][1] ), 
	.D(n236), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[6][0]  (.SI(\memory[5][7] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[6][0] ), 
	.D(n235), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \memory_reg[12][7]  (.SI(\memory[12][6] ), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[12][7] ), 
	.D(n290), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[12][6]  (.SI(\memory[12][5] ), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[12][6] ), 
	.D(n289), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[12][5]  (.SI(\memory[12][4] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[12][5] ), 
	.D(n288), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[12][4]  (.SI(\memory[12][3] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[12][4] ), 
	.D(n287), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[12][3]  (.SI(\memory[12][2] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[12][3] ), 
	.D(n286), 
	.CK(REF_CLK_M__L5_N8));
   SDFFRQX2M \memory_reg[12][2]  (.SI(\memory[12][1] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[12][2] ), 
	.D(n285), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[12][1]  (.SI(\memory[12][0] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[12][1] ), 
	.D(n284), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[12][0]  (.SI(\memory[11][7] ), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[12][0] ), 
	.D(n283), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[8][7]  (.SI(test_si2), 
	.SE(n373), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(\memory[8][7] ), 
	.D(n258), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[8][6]  (.SI(\memory[8][5] ), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[8][6] ), 
	.D(n257), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[8][5]  (.SI(\memory[8][4] ), 
	.SE(n371), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[8][5] ), 
	.D(n256), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[8][4]  (.SI(\memory[8][3] ), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[8][4] ), 
	.D(n255), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[8][3]  (.SI(\memory[8][2] ), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[8][3] ), 
	.D(n254), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[8][2]  (.SI(\memory[8][1] ), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(\memory[8][2] ), 
	.D(n253), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[8][1]  (.SI(\memory[8][0] ), 
	.SE(n371), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(\memory[8][1] ), 
	.D(n252), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[8][0]  (.SI(\memory[7][7] ), 
	.SE(n370), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(\memory[8][0] ), 
	.D(n251), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[4][7]  (.SI(\memory[4][6] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[4][7] ), 
	.D(n226), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[4][6]  (.SI(\memory[4][5] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[4][6] ), 
	.D(n225), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[4][5]  (.SI(\memory[4][4] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[4][5] ), 
	.D(n224), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[4][4]  (.SI(\memory[4][3] ), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[4][4] ), 
	.D(n223), 
	.CK(REF_CLK_M__L5_N12));
   SDFFRQX2M \memory_reg[4][3]  (.SI(\memory[4][2] ), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[4][3] ), 
	.D(n222), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[4][2]  (.SI(\memory[4][1] ), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[4][2] ), 
	.D(n221), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[4][1]  (.SI(\memory[4][0] ), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[4][1] ), 
	.D(n220), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[4][0]  (.SI(REG3[7]), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(\memory[4][0] ), 
	.D(n219), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \RdData_reg[7]  (.SI(RdData[6]), 
	.SE(n373), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(RdData[7]), 
	.D(n185), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \RdData_reg[6]  (.SI(RdData[5]), 
	.SE(n372), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(RdData[6]), 
	.D(n184), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \RdData_reg[5]  (.SI(RdData[4]), 
	.SE(n371), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(RdData[5]), 
	.D(n183), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \RdData_reg[4]  (.SI(RdData[3]), 
	.SE(n370), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(RdData[4]), 
	.D(n182), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \RdData_reg[3]  (.SI(RdData[2]), 
	.SE(n373), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(RdData[3]), 
	.D(n181), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \RdData_reg[2]  (.SI(RdData[1]), 
	.SE(n372), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(RdData[2]), 
	.D(n180), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \RdData_reg[1]  (.SI(RdData[0]), 
	.SE(n371), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(RdData[1]), 
	.D(n179), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \RdData_reg[0]  (.SI(RdData_VLD), 
	.SE(n370), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(RdData[0]), 
	.D(n178), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M RdData_VLD_reg (.SI(test_si1), 
	.SE(n373), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(RdData_VLD), 
	.D(n186), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \memory_reg[3][0]  (.SI(REG2[7]), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG3[0]), 
	.D(n211), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \memory_reg[2][0]  (.SI(REG1[7]), 
	.SE(n371), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(REG2[0]), 
	.D(n203), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \memory_reg[2][1]  (.SI(REG2[0]), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG2[1]), 
	.D(n204), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \memory_reg[1][7]  (.SI(REG1[6]), 
	.SE(n373), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(REG1[7]), 
	.D(n202), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[1][6]  (.SI(REG1[5]), 
	.SE(n372), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(REG1[6]), 
	.D(n201), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[1][1]  (.SI(REG1[0]), 
	.SE(n371), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG1[1]), 
	.D(n196), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[0][7]  (.SI(REG0[6]), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG0[7]), 
	.D(n194), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[0][6]  (.SI(REG0[5]), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG0[6]), 
	.D(n193), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[0][5]  (.SI(REG0[4]), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG0[5]), 
	.D(n192), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[0][4]  (.SI(REG0[3]), 
	.SE(n371), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG0[4]), 
	.D(n191), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[0][3]  (.SI(REG0[2]), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG0[3]), 
	.D(n190), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[0][2]  (.SI(REG0[1]), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG0[2]), 
	.D(n189), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[0][1]  (.SI(REG0[0]), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG0[1]), 
	.D(n188), 
	.CK(CLK));
   SDFFRQX2M \memory_reg[0][0]  (.SI(RdData[7]), 
	.SE(n371), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(REG0[0]), 
	.D(n187), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[1][4]  (.SI(REG1[3]), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG1[4]), 
	.D(n199), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[1][5]  (.SI(REG1[4]), 
	.SE(n373), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG1[5]), 
	.D(n200), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[3][7]  (.SI(REG3[6]), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG3[7]), 
	.D(n218), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \memory_reg[3][6]  (.SI(REG3[5]), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG3[6]), 
	.D(n217), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \memory_reg[3][2]  (.SI(REG3[1]), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG3[2]), 
	.D(n213), 
	.CK(REF_CLK_M__L5_N15));
   SDFFRQX2M \memory_reg[3][3]  (.SI(REG3[2]), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG3[3]), 
	.D(n214), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \memory_reg[3][4]  (.SI(REG3[3]), 
	.SE(n372), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG3[4]), 
	.D(n215), 
	.CK(REF_CLK_M__L5_N3));
   SDFFSQX2M \memory_reg[3][5]  (.SN(FE_OFN2_M_Domain1_SYNC_RST), 
	.SI(REG3[4]), 
	.SE(test_se), 
	.Q(REG3[5]), 
	.D(n216), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \memory_reg[3][1]  (.SI(REG3[0]), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG3[1]), 
	.D(n212), 
	.CK(REF_CLK_M__L5_N14));
   SDFFSQX2M \memory_reg[2][7]  (.SN(FE_OFN2_M_Domain1_SYNC_RST), 
	.SI(REG2[6]), 
	.SE(n370), 
	.Q(REG2[7]), 
	.D(n210), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \memory_reg[2][3]  (.SI(REG2[2]), 
	.SE(n370), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG2[3]), 
	.D(n206), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \memory_reg[2][4]  (.SI(REG2[3]), 
	.SE(n373), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG2[4]), 
	.D(n207), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \memory_reg[2][2]  (.SI(REG2[1]), 
	.SE(n372), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(REG2[2]), 
	.D(n205), 
	.CK(REF_CLK_M__L5_N14));
   SDFFRQX2M \memory_reg[2][6]  (.SI(REG2[5]), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG2[6]), 
	.D(n209), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \memory_reg[1][2]  (.SI(REG1[1]), 
	.SE(n370), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG1[2]), 
	.D(n197), 
	.CK(REF_CLK_M__L5_N9));
   SDFFRQX2M \memory_reg[1][3]  (.SI(REG1[2]), 
	.SE(n373), 
	.RN(FE_OFN4_M_Domain1_SYNC_RST), 
	.Q(REG1[3]), 
	.D(n198), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[1][0]  (.SI(REG0[7]), 
	.SE(n372), 
	.RN(FE_OFN3_M_Domain1_SYNC_RST), 
	.Q(REG1[0]), 
	.D(n195), 
	.CK(REF_CLK_M__L5_N13));
   SDFFRQX2M \memory_reg[2][5]  (.SI(REG2[4]), 
	.SE(n371), 
	.RN(FE_OFN2_M_Domain1_SYNC_RST), 
	.Q(REG2[5]), 
	.D(n208), 
	.CK(REF_CLK_M__L5_N3));
   NOR2X2M U140 (.Y(n155), 
	.B(N13), 
	.A(n341));
   NOR2X2M U141 (.Y(n153), 
	.B(N13), 
	.A(N12));
   INVX4M U142 (.Y(n338), 
	.A(n340));
   INVX2M U143 (.Y(n336), 
	.A(n341));
   INVX4M U144 (.Y(n339), 
	.A(n340));
   NAND2X2M U147 (.Y(n173), 
	.B(n159), 
	.A(n168));
   NAND2X2M U148 (.Y(n174), 
	.B(n159), 
	.A(n170));
   NAND2X2M U149 (.Y(n175), 
	.B(n162), 
	.A(n168));
   NAND2X2M U150 (.Y(n177), 
	.B(n162), 
	.A(n170));
   NAND2X2M U151 (.Y(n154), 
	.B(n156), 
	.A(n155));
   NAND2X2M U152 (.Y(n157), 
	.B(n152), 
	.A(n155));
   NAND2X2M U153 (.Y(n158), 
	.B(n156), 
	.A(n159));
   NAND2X2M U154 (.Y(n160), 
	.B(n152), 
	.A(n159));
   NAND2X2M U155 (.Y(n161), 
	.B(n156), 
	.A(n162));
   NAND2X2M U156 (.Y(n163), 
	.B(n152), 
	.A(n162));
   NAND2X2M U157 (.Y(n167), 
	.B(n153), 
	.A(n168));
   NAND2X2M U158 (.Y(n169), 
	.B(n153), 
	.A(n170));
   NAND2X2M U159 (.Y(n171), 
	.B(n155), 
	.A(n168));
   NAND2X2M U160 (.Y(n172), 
	.B(n155), 
	.A(n170));
   NAND2X2M U161 (.Y(n151), 
	.B(n153), 
	.A(n152));
   NAND2X2M U162 (.Y(n150), 
	.B(n156), 
	.A(n153));
   AND2X2M U163 (.Y(n152), 
	.B(N11), 
	.A(n164));
   AND2X2M U164 (.Y(n170), 
	.B(N11), 
	.A(n176));
   INVX2M U165 (.Y(n365), 
	.A(n165));
   NAND2X2M U176 (.Y(n165), 
	.B(n366), 
	.A(RdEn));
   NOR2X2M U177 (.Y(n166), 
	.B(RdEn), 
	.A(n366));
   AND2X2M U178 (.Y(n159), 
	.B(n341), 
	.A(N13));
   AND2X2M U179 (.Y(n162), 
	.B(N12), 
	.A(N13));
   AND2X2M U180 (.Y(n156), 
	.B(n340), 
	.A(n164));
   NOR2BX2M U181 (.Y(n176), 
	.B(N14), 
	.AN(n166));
   AND2X2M U182 (.Y(n168), 
	.B(n340), 
	.A(n176));
   AND2X2M U183 (.Y(n164), 
	.B(n166), 
	.A(N14));
   INVX2M U184 (.Y(n366), 
	.A(WrEn));
   AO22X1M U190 (.Y(n178), 
	.B1(n165), 
	.B0(RdData[0]), 
	.A1(n365), 
	.A0(N43));
   MX4X1M U191 (.Y(N43), 
	.S1(N13), 
	.S0(N14), 
	.D(n138), 
	.C(n140), 
	.B(n139), 
	.A(n141));
   MX4X1M U192 (.Y(n141), 
	.S1(N12), 
	.S0(N11), 
	.D(REG3[0]), 
	.C(REG2[0]), 
	.B(REG1[0]), 
	.A(REG0[0]));
   MX4X1M U193 (.Y(n139), 
	.S1(N12), 
	.S0(N11), 
	.D(\memory[11][0] ), 
	.C(\memory[10][0] ), 
	.B(\memory[9][0] ), 
	.A(\memory[8][0] ));
   AO22X1M U194 (.Y(n179), 
	.B1(n165), 
	.B0(RdData[1]), 
	.A1(n365), 
	.A0(N42));
   MX4X1M U195 (.Y(N42), 
	.S1(N13), 
	.S0(N14), 
	.D(n142), 
	.C(n144), 
	.B(n143), 
	.A(n145));
   MX4X1M U196 (.Y(n143), 
	.S1(N12), 
	.S0(N11), 
	.D(\memory[11][1] ), 
	.C(\memory[10][1] ), 
	.B(\memory[9][1] ), 
	.A(\memory[8][1] ));
   MX4X1M U197 (.Y(n142), 
	.S1(n336), 
	.S0(n338), 
	.D(\memory[15][1] ), 
	.C(\memory[14][1] ), 
	.B(\memory[13][1] ), 
	.A(\memory[12][1] ));
   AO22X1M U198 (.Y(n180), 
	.B1(n165), 
	.B0(RdData[2]), 
	.A1(n365), 
	.A0(N41));
   MX4X1M U199 (.Y(N41), 
	.S1(N13), 
	.S0(N14), 
	.D(n146), 
	.C(n148), 
	.B(n147), 
	.A(n149));
   MX4X1M U200 (.Y(n149), 
	.S1(n336), 
	.S0(n338), 
	.D(REG3[2]), 
	.C(REG2[2]), 
	.B(REG1[2]), 
	.A(REG0[2]));
   MX4X1M U201 (.Y(n147), 
	.S1(n336), 
	.S0(n338), 
	.D(\memory[11][2] ), 
	.C(\memory[10][2] ), 
	.B(\memory[9][2] ), 
	.A(\memory[8][2] ));
   AO22X1M U202 (.Y(n181), 
	.B1(n165), 
	.B0(RdData[3]), 
	.A1(n365), 
	.A0(N40));
   MX4X1M U203 (.Y(N40), 
	.S1(N13), 
	.S0(N14), 
	.D(n315), 
	.C(n317), 
	.B(n316), 
	.A(n318));
   MX4X1M U204 (.Y(n318), 
	.S1(n336), 
	.S0(n338), 
	.D(REG3[3]), 
	.C(REG2[3]), 
	.B(REG1[3]), 
	.A(REG0[3]));
   MX4X1M U205 (.Y(n316), 
	.S1(n336), 
	.S0(n338), 
	.D(\memory[11][3] ), 
	.C(\memory[10][3] ), 
	.B(\memory[9][3] ), 
	.A(\memory[8][3] ));
   AO22X1M U206 (.Y(n182), 
	.B1(n165), 
	.B0(RdData[4]), 
	.A1(n365), 
	.A0(N39));
   MX4X1M U207 (.Y(N39), 
	.S1(N13), 
	.S0(N14), 
	.D(n319), 
	.C(n321), 
	.B(n320), 
	.A(n322));
   MX4X1M U208 (.Y(n322), 
	.S1(n336), 
	.S0(n339), 
	.D(REG3[4]), 
	.C(REG2[4]), 
	.B(REG1[4]), 
	.A(REG0[4]));
   MX4X1M U209 (.Y(n320), 
	.S1(n336), 
	.S0(n338), 
	.D(\memory[11][4] ), 
	.C(\memory[10][4] ), 
	.B(\memory[9][4] ), 
	.A(\memory[8][4] ));
   AO22X1M U210 (.Y(n183), 
	.B1(n165), 
	.B0(RdData[5]), 
	.A1(n365), 
	.A0(N38));
   MX4X1M U211 (.Y(N38), 
	.S1(N13), 
	.S0(N14), 
	.D(n323), 
	.C(n325), 
	.B(n324), 
	.A(n326));
   MX4X1M U212 (.Y(n326), 
	.S1(N12), 
	.S0(n339), 
	.D(REG3[5]), 
	.C(REG2[5]), 
	.B(REG1[5]), 
	.A(REG0[5]));
   MX4X1M U213 (.Y(n324), 
	.S1(N12), 
	.S0(n339), 
	.D(\memory[11][5] ), 
	.C(\memory[10][5] ), 
	.B(\memory[9][5] ), 
	.A(\memory[8][5] ));
   AO22X1M U214 (.Y(n184), 
	.B1(n165), 
	.B0(RdData[6]), 
	.A1(n365), 
	.A0(N37));
   MX4X1M U215 (.Y(N37), 
	.S1(N13), 
	.S0(N14), 
	.D(n327), 
	.C(n329), 
	.B(n328), 
	.A(n330));
   MX4X1M U216 (.Y(n330), 
	.S1(N12), 
	.S0(n339), 
	.D(REG3[6]), 
	.C(REG2[6]), 
	.B(REG1[6]), 
	.A(REG0[6]));
   MX4X1M U217 (.Y(n328), 
	.S1(N12), 
	.S0(n339), 
	.D(\memory[11][6] ), 
	.C(\memory[10][6] ), 
	.B(\memory[9][6] ), 
	.A(\memory[8][6] ));
   AO22X1M U218 (.Y(n185), 
	.B1(n165), 
	.B0(RdData[7]), 
	.A1(n365), 
	.A0(N36));
   MX4X1M U219 (.Y(N36), 
	.S1(N13), 
	.S0(N14), 
	.D(n331), 
	.C(n333), 
	.B(n332), 
	.A(n334));
   MX4X1M U220 (.Y(n334), 
	.S1(N12), 
	.S0(n339), 
	.D(REG3[7]), 
	.C(REG2[7]), 
	.B(REG1[7]), 
	.A(REG0[7]));
   MX4X1M U221 (.Y(n332), 
	.S1(N12), 
	.S0(n339), 
	.D(\memory[11][7] ), 
	.C(\memory[10][7] ), 
	.B(\memory[9][7] ), 
	.A(\memory[8][7] ));
   MX4X1M U222 (.Y(n145), 
	.S1(N12), 
	.S0(n338), 
	.D(REG3[1]), 
	.C(REG2[1]), 
	.B(REG1[1]), 
	.A(REG0[1]));
   MX4X1M U223 (.Y(n140), 
	.S1(N12), 
	.S0(N11), 
	.D(\memory[7][0] ), 
	.C(\memory[6][0] ), 
	.B(\memory[5][0] ), 
	.A(\memory[4][0] ));
   MX4X1M U224 (.Y(n144), 
	.S1(N12), 
	.S0(n338), 
	.D(\memory[7][1] ), 
	.C(\memory[6][1] ), 
	.B(\memory[5][1] ), 
	.A(\memory[4][1] ));
   MX4X1M U225 (.Y(n148), 
	.S1(n336), 
	.S0(n338), 
	.D(\memory[7][2] ), 
	.C(\memory[6][2] ), 
	.B(\memory[5][2] ), 
	.A(\memory[4][2] ));
   MX4X1M U226 (.Y(n317), 
	.S1(n336), 
	.S0(n338), 
	.D(\memory[7][3] ), 
	.C(\memory[6][3] ), 
	.B(\memory[5][3] ), 
	.A(\memory[4][3] ));
   MX4X1M U227 (.Y(n321), 
	.S1(n336), 
	.S0(n338), 
	.D(\memory[7][4] ), 
	.C(\memory[6][4] ), 
	.B(\memory[5][4] ), 
	.A(\memory[4][4] ));
   MX4X1M U228 (.Y(n325), 
	.S1(N12), 
	.S0(n339), 
	.D(\memory[7][5] ), 
	.C(\memory[6][5] ), 
	.B(\memory[5][5] ), 
	.A(\memory[4][5] ));
   MX4X1M U229 (.Y(n329), 
	.S1(N12), 
	.S0(n339), 
	.D(\memory[7][6] ), 
	.C(\memory[6][6] ), 
	.B(\memory[5][6] ), 
	.A(\memory[4][6] ));
   MX4X1M U230 (.Y(n333), 
	.S1(N12), 
	.S0(n339), 
	.D(\memory[7][7] ), 
	.C(\memory[6][7] ), 
	.B(\memory[5][7] ), 
	.A(\memory[4][7] ));
   MX4X1M U231 (.Y(n138), 
	.S1(n336), 
	.S0(n339), 
	.D(\memory[15][0] ), 
	.C(\memory[14][0] ), 
	.B(\memory[13][0] ), 
	.A(\memory[12][0] ));
   MX4X1M U232 (.Y(n146), 
	.S1(n336), 
	.S0(n338), 
	.D(\memory[15][2] ), 
	.C(\memory[14][2] ), 
	.B(\memory[13][2] ), 
	.A(\memory[12][2] ));
   MX4X1M U233 (.Y(n315), 
	.S1(n336), 
	.S0(n338), 
	.D(\memory[15][3] ), 
	.C(\memory[14][3] ), 
	.B(\memory[13][3] ), 
	.A(\memory[12][3] ));
   MX4X1M U234 (.Y(n319), 
	.S1(n336), 
	.S0(n338), 
	.D(\memory[15][4] ), 
	.C(\memory[14][4] ), 
	.B(\memory[13][4] ), 
	.A(\memory[12][4] ));
   MX4X1M U235 (.Y(n323), 
	.S1(N12), 
	.S0(n339), 
	.D(\memory[15][5] ), 
	.C(\memory[14][5] ), 
	.B(\memory[13][5] ), 
	.A(\memory[12][5] ));
   MX4X1M U236 (.Y(n327), 
	.S1(N12), 
	.S0(n339), 
	.D(\memory[15][6] ), 
	.C(\memory[14][6] ), 
	.B(\memory[13][6] ), 
	.A(\memory[12][6] ));
   MX4X1M U237 (.Y(n331), 
	.S1(N12), 
	.S0(n339), 
	.D(\memory[15][7] ), 
	.C(\memory[14][7] ), 
	.B(\memory[13][7] ), 
	.A(\memory[12][7] ));
   INVX2M U238 (.Y(n340), 
	.A(N11));
   INVX2M U239 (.Y(n363), 
	.A(WrData[1]));
   INVX2M U240 (.Y(n362), 
	.A(WrData[2]));
   INVX2M U241 (.Y(n361), 
	.A(WrData[3]));
   INVX2M U242 (.Y(n364), 
	.A(WrData[0]));
   INVX2M U243 (.Y(n360), 
	.A(WrData[4]));
   INVX2M U244 (.Y(n359), 
	.A(WrData[5]));
   INVX2M U245 (.Y(n358), 
	.A(WrData[6]));
   INVX2M U246 (.Y(n357), 
	.A(WrData[7]));
   OAI2BB2X1M U247 (.Y(n251), 
	.B1(n364), 
	.B0(n150), 
	.A1N(n150), 
	.A0N(\memory[8][0] ));
   OAI2BB2X1M U248 (.Y(n252), 
	.B1(n363), 
	.B0(n150), 
	.A1N(n150), 
	.A0N(\memory[8][1] ));
   OAI2BB2X1M U249 (.Y(n253), 
	.B1(n362), 
	.B0(n150), 
	.A1N(n150), 
	.A0N(\memory[8][2] ));
   OAI2BB2X1M U250 (.Y(n254), 
	.B1(n361), 
	.B0(n150), 
	.A1N(n150), 
	.A0N(\memory[8][3] ));
   OAI2BB2X1M U251 (.Y(n255), 
	.B1(n360), 
	.B0(n150), 
	.A1N(n150), 
	.A0N(\memory[8][4] ));
   OAI2BB2X1M U252 (.Y(n256), 
	.B1(n359), 
	.B0(n150), 
	.A1N(n150), 
	.A0N(\memory[8][5] ));
   OAI2BB2X1M U253 (.Y(n257), 
	.B1(n358), 
	.B0(n150), 
	.A1N(n150), 
	.A0N(\memory[8][6] ));
   OAI2BB2X1M U254 (.Y(n258), 
	.B1(n357), 
	.B0(n150), 
	.A1N(n150), 
	.A0N(\memory[8][7] ));
   OAI2BB2X1M U255 (.Y(n267), 
	.B1(n154), 
	.B0(n364), 
	.A1N(n154), 
	.A0N(\memory[10][0] ));
   OAI2BB2X1M U256 (.Y(n268), 
	.B1(n154), 
	.B0(n363), 
	.A1N(n154), 
	.A0N(\memory[10][1] ));
   OAI2BB2X1M U257 (.Y(n269), 
	.B1(n154), 
	.B0(n362), 
	.A1N(n154), 
	.A0N(\memory[10][2] ));
   OAI2BB2X1M U258 (.Y(n270), 
	.B1(n154), 
	.B0(n361), 
	.A1N(n154), 
	.A0N(\memory[10][3] ));
   OAI2BB2X1M U259 (.Y(n271), 
	.B1(n154), 
	.B0(n360), 
	.A1N(n154), 
	.A0N(\memory[10][4] ));
   OAI2BB2X1M U260 (.Y(n272), 
	.B1(n154), 
	.B0(n359), 
	.A1N(n154), 
	.A0N(\memory[10][5] ));
   OAI2BB2X1M U261 (.Y(n273), 
	.B1(n154), 
	.B0(n358), 
	.A1N(n154), 
	.A0N(\memory[10][6] ));
   OAI2BB2X1M U262 (.Y(n274), 
	.B1(n154), 
	.B0(n357), 
	.A1N(n154), 
	.A0N(\memory[10][7] ));
   OAI2BB2X1M U263 (.Y(n275), 
	.B1(n157), 
	.B0(n364), 
	.A1N(n157), 
	.A0N(\memory[11][0] ));
   OAI2BB2X1M U264 (.Y(n276), 
	.B1(n157), 
	.B0(n363), 
	.A1N(n157), 
	.A0N(\memory[11][1] ));
   OAI2BB2X1M U265 (.Y(n277), 
	.B1(n157), 
	.B0(n362), 
	.A1N(n157), 
	.A0N(\memory[11][2] ));
   OAI2BB2X1M U266 (.Y(n278), 
	.B1(n157), 
	.B0(n361), 
	.A1N(n157), 
	.A0N(\memory[11][3] ));
   OAI2BB2X1M U267 (.Y(n279), 
	.B1(n157), 
	.B0(n360), 
	.A1N(n157), 
	.A0N(\memory[11][4] ));
   OAI2BB2X1M U268 (.Y(n280), 
	.B1(n157), 
	.B0(n359), 
	.A1N(n157), 
	.A0N(\memory[11][5] ));
   OAI2BB2X1M U269 (.Y(n281), 
	.B1(n157), 
	.B0(n358), 
	.A1N(n157), 
	.A0N(\memory[11][6] ));
   OAI2BB2X1M U270 (.Y(n282), 
	.B1(n157), 
	.B0(n357), 
	.A1N(n157), 
	.A0N(\memory[11][7] ));
   OAI2BB2X1M U271 (.Y(n259), 
	.B1(n364), 
	.B0(n151), 
	.A1N(n151), 
	.A0N(\memory[9][0] ));
   OAI2BB2X1M U272 (.Y(n260), 
	.B1(n363), 
	.B0(n151), 
	.A1N(n151), 
	.A0N(\memory[9][1] ));
   OAI2BB2X1M U273 (.Y(n261), 
	.B1(n362), 
	.B0(n151), 
	.A1N(n151), 
	.A0N(\memory[9][2] ));
   OAI2BB2X1M U274 (.Y(n262), 
	.B1(n361), 
	.B0(n151), 
	.A1N(n151), 
	.A0N(\memory[9][3] ));
   OAI2BB2X1M U275 (.Y(n263), 
	.B1(n360), 
	.B0(n151), 
	.A1N(n151), 
	.A0N(\memory[9][4] ));
   OAI2BB2X1M U276 (.Y(n264), 
	.B1(n359), 
	.B0(n151), 
	.A1N(n151), 
	.A0N(\memory[9][5] ));
   OAI2BB2X1M U277 (.Y(n265), 
	.B1(n358), 
	.B0(n151), 
	.A1N(n151), 
	.A0N(\memory[9][6] ));
   OAI2BB2X1M U278 (.Y(n187), 
	.B1(n167), 
	.B0(n364), 
	.A1N(n167), 
	.A0N(REG0[0]));
   OAI2BB2X1M U279 (.Y(n188), 
	.B1(n167), 
	.B0(n363), 
	.A1N(n167), 
	.A0N(REG0[1]));
   OAI2BB2X1M U280 (.Y(n189), 
	.B1(n167), 
	.B0(n362), 
	.A1N(n167), 
	.A0N(REG0[2]));
   OAI2BB2X1M U281 (.Y(n190), 
	.B1(n167), 
	.B0(n361), 
	.A1N(n167), 
	.A0N(REG0[3]));
   OAI2BB2X1M U282 (.Y(n191), 
	.B1(n167), 
	.B0(n360), 
	.A1N(n167), 
	.A0N(REG0[4]));
   OAI2BB2X1M U283 (.Y(n192), 
	.B1(n167), 
	.B0(n359), 
	.A1N(n167), 
	.A0N(REG0[5]));
   OAI2BB2X1M U284 (.Y(n193), 
	.B1(n167), 
	.B0(n358), 
	.A1N(n167), 
	.A0N(REG0[6]));
   OAI2BB2X1M U285 (.Y(n194), 
	.B1(n167), 
	.B0(n357), 
	.A1N(n167), 
	.A0N(REG0[7]));
   OAI2BB2X1M U286 (.Y(n195), 
	.B1(n169), 
	.B0(n364), 
	.A1N(n169), 
	.A0N(REG1[0]));
   OAI2BB2X1M U287 (.Y(n196), 
	.B1(n169), 
	.B0(n363), 
	.A1N(n169), 
	.A0N(REG1[1]));
   OAI2BB2X1M U288 (.Y(n197), 
	.B1(n169), 
	.B0(n362), 
	.A1N(n169), 
	.A0N(REG1[2]));
   OAI2BB2X1M U289 (.Y(n198), 
	.B1(n169), 
	.B0(n361), 
	.A1N(n169), 
	.A0N(REG1[3]));
   OAI2BB2X1M U290 (.Y(n199), 
	.B1(n169), 
	.B0(n360), 
	.A1N(n169), 
	.A0N(REG1[4]));
   OAI2BB2X1M U291 (.Y(n200), 
	.B1(n169), 
	.B0(n359), 
	.A1N(n169), 
	.A0N(REG1[5]));
   OAI2BB2X1M U292 (.Y(n201), 
	.B1(n169), 
	.B0(n358), 
	.A1N(n169), 
	.A0N(REG1[6]));
   OAI2BB2X1M U293 (.Y(n202), 
	.B1(n169), 
	.B0(n357), 
	.A1N(n169), 
	.A0N(REG1[7]));
   OAI2BB2X1M U294 (.Y(n203), 
	.B1(n171), 
	.B0(n364), 
	.A1N(n171), 
	.A0N(REG2[0]));
   OAI2BB2X1M U295 (.Y(n204), 
	.B1(n171), 
	.B0(n363), 
	.A1N(n171), 
	.A0N(REG2[1]));
   OAI2BB2X1M U296 (.Y(n205), 
	.B1(n171), 
	.B0(n362), 
	.A1N(n171), 
	.A0N(REG2[2]));
   OAI2BB2X1M U297 (.Y(n206), 
	.B1(n171), 
	.B0(n361), 
	.A1N(n171), 
	.A0N(REG2[3]));
   OAI2BB2X1M U298 (.Y(n207), 
	.B1(n171), 
	.B0(n360), 
	.A1N(n171), 
	.A0N(REG2[4]));
   OAI2BB2X1M U299 (.Y(n208), 
	.B1(n171), 
	.B0(n359), 
	.A1N(n171), 
	.A0N(REG2[5]));
   OAI2BB2X1M U300 (.Y(n209), 
	.B1(n171), 
	.B0(n358), 
	.A1N(n171), 
	.A0N(REG2[6]));
   OAI2BB2X1M U301 (.Y(n211), 
	.B1(n172), 
	.B0(n364), 
	.A1N(n172), 
	.A0N(REG3[0]));
   OAI2BB2X1M U302 (.Y(n212), 
	.B1(n172), 
	.B0(n363), 
	.A1N(n172), 
	.A0N(REG3[1]));
   OAI2BB2X1M U303 (.Y(n213), 
	.B1(n172), 
	.B0(n362), 
	.A1N(n172), 
	.A0N(REG3[2]));
   OAI2BB2X1M U304 (.Y(n214), 
	.B1(n172), 
	.B0(n361), 
	.A1N(n172), 
	.A0N(REG3[3]));
   OAI2BB2X1M U305 (.Y(n215), 
	.B1(n172), 
	.B0(n360), 
	.A1N(n172), 
	.A0N(REG3[4]));
   OAI2BB2X1M U306 (.Y(n217), 
	.B1(n172), 
	.B0(n358), 
	.A1N(n172), 
	.A0N(REG3[6]));
   OAI2BB2X1M U307 (.Y(n218), 
	.B1(n172), 
	.B0(n357), 
	.A1N(n172), 
	.A0N(REG3[7]));
   OAI2BB2X1M U308 (.Y(n266), 
	.B1(n151), 
	.B0(n357), 
	.A1N(n151), 
	.A0N(\memory[9][7] ));
   OAI2BB2X1M U309 (.Y(n210), 
	.B1(n171), 
	.B0(n357), 
	.A1N(n171), 
	.A0N(REG2[7]));
   OAI2BB2X1M U310 (.Y(n216), 
	.B1(n172), 
	.B0(n359), 
	.A1N(n172), 
	.A0N(REG3[5]));
   OAI2BB2X1M U311 (.Y(n219), 
	.B1(n173), 
	.B0(n364), 
	.A1N(n173), 
	.A0N(\memory[4][0] ));
   OAI2BB2X1M U312 (.Y(n220), 
	.B1(n173), 
	.B0(n363), 
	.A1N(n173), 
	.A0N(\memory[4][1] ));
   OAI2BB2X1M U313 (.Y(n221), 
	.B1(n173), 
	.B0(n362), 
	.A1N(n173), 
	.A0N(\memory[4][2] ));
   OAI2BB2X1M U314 (.Y(n222), 
	.B1(n173), 
	.B0(n361), 
	.A1N(n173), 
	.A0N(\memory[4][3] ));
   OAI2BB2X1M U315 (.Y(n223), 
	.B1(n173), 
	.B0(n360), 
	.A1N(n173), 
	.A0N(\memory[4][4] ));
   OAI2BB2X1M U316 (.Y(n224), 
	.B1(n173), 
	.B0(n359), 
	.A1N(n173), 
	.A0N(\memory[4][5] ));
   OAI2BB2X1M U317 (.Y(n225), 
	.B1(n173), 
	.B0(n358), 
	.A1N(n173), 
	.A0N(\memory[4][6] ));
   OAI2BB2X1M U318 (.Y(n226), 
	.B1(n173), 
	.B0(n357), 
	.A1N(n173), 
	.A0N(\memory[4][7] ));
   OAI2BB2X1M U319 (.Y(n227), 
	.B1(n174), 
	.B0(n364), 
	.A1N(n174), 
	.A0N(\memory[5][0] ));
   OAI2BB2X1M U320 (.Y(n228), 
	.B1(n174), 
	.B0(n363), 
	.A1N(n174), 
	.A0N(\memory[5][1] ));
   OAI2BB2X1M U321 (.Y(n229), 
	.B1(n174), 
	.B0(n362), 
	.A1N(n174), 
	.A0N(\memory[5][2] ));
   OAI2BB2X1M U322 (.Y(n230), 
	.B1(n174), 
	.B0(n361), 
	.A1N(n174), 
	.A0N(\memory[5][3] ));
   OAI2BB2X1M U323 (.Y(n231), 
	.B1(n174), 
	.B0(n360), 
	.A1N(n174), 
	.A0N(\memory[5][4] ));
   OAI2BB2X1M U324 (.Y(n232), 
	.B1(n174), 
	.B0(n359), 
	.A1N(n174), 
	.A0N(\memory[5][5] ));
   OAI2BB2X1M U325 (.Y(n233), 
	.B1(n174), 
	.B0(n358), 
	.A1N(n174), 
	.A0N(\memory[5][6] ));
   OAI2BB2X1M U326 (.Y(n234), 
	.B1(n174), 
	.B0(n357), 
	.A1N(n174), 
	.A0N(\memory[5][7] ));
   OAI2BB2X1M U327 (.Y(n235), 
	.B1(n175), 
	.B0(n364), 
	.A1N(n175), 
	.A0N(\memory[6][0] ));
   OAI2BB2X1M U328 (.Y(n236), 
	.B1(n175), 
	.B0(n363), 
	.A1N(n175), 
	.A0N(\memory[6][1] ));
   OAI2BB2X1M U329 (.Y(n237), 
	.B1(n175), 
	.B0(n362), 
	.A1N(n175), 
	.A0N(\memory[6][2] ));
   OAI2BB2X1M U330 (.Y(n238), 
	.B1(n175), 
	.B0(n361), 
	.A1N(n175), 
	.A0N(\memory[6][3] ));
   OAI2BB2X1M U331 (.Y(n239), 
	.B1(n175), 
	.B0(n360), 
	.A1N(n175), 
	.A0N(\memory[6][4] ));
   OAI2BB2X1M U332 (.Y(n240), 
	.B1(n175), 
	.B0(n359), 
	.A1N(n175), 
	.A0N(\memory[6][5] ));
   OAI2BB2X1M U333 (.Y(n241), 
	.B1(n175), 
	.B0(n358), 
	.A1N(n175), 
	.A0N(\memory[6][6] ));
   OAI2BB2X1M U334 (.Y(n242), 
	.B1(n175), 
	.B0(n357), 
	.A1N(n175), 
	.A0N(\memory[6][7] ));
   OAI2BB2X1M U335 (.Y(n243), 
	.B1(n177), 
	.B0(n364), 
	.A1N(n177), 
	.A0N(\memory[7][0] ));
   OAI2BB2X1M U336 (.Y(n244), 
	.B1(n177), 
	.B0(n363), 
	.A1N(n177), 
	.A0N(\memory[7][1] ));
   OAI2BB2X1M U337 (.Y(n245), 
	.B1(n177), 
	.B0(n362), 
	.A1N(n177), 
	.A0N(\memory[7][2] ));
   OAI2BB2X1M U338 (.Y(n246), 
	.B1(n177), 
	.B0(n361), 
	.A1N(n177), 
	.A0N(\memory[7][3] ));
   OAI2BB2X1M U339 (.Y(n247), 
	.B1(n177), 
	.B0(n360), 
	.A1N(n177), 
	.A0N(\memory[7][4] ));
   OAI2BB2X1M U340 (.Y(n248), 
	.B1(n177), 
	.B0(n359), 
	.A1N(n177), 
	.A0N(\memory[7][5] ));
   OAI2BB2X1M U341 (.Y(n249), 
	.B1(n177), 
	.B0(n358), 
	.A1N(n177), 
	.A0N(\memory[7][6] ));
   OAI2BB2X1M U342 (.Y(n250), 
	.B1(n177), 
	.B0(n357), 
	.A1N(n177), 
	.A0N(\memory[7][7] ));
   OAI2BB2X1M U343 (.Y(n283), 
	.B1(n158), 
	.B0(n364), 
	.A1N(n158), 
	.A0N(\memory[12][0] ));
   OAI2BB2X1M U344 (.Y(n284), 
	.B1(n158), 
	.B0(n363), 
	.A1N(n158), 
	.A0N(\memory[12][1] ));
   OAI2BB2X1M U345 (.Y(n285), 
	.B1(n158), 
	.B0(n362), 
	.A1N(n158), 
	.A0N(\memory[12][2] ));
   OAI2BB2X1M U346 (.Y(n286), 
	.B1(n158), 
	.B0(n361), 
	.A1N(n158), 
	.A0N(\memory[12][3] ));
   OAI2BB2X1M U347 (.Y(n287), 
	.B1(n158), 
	.B0(n360), 
	.A1N(n158), 
	.A0N(\memory[12][4] ));
   OAI2BB2X1M U348 (.Y(n288), 
	.B1(n158), 
	.B0(n359), 
	.A1N(n158), 
	.A0N(\memory[12][5] ));
   OAI2BB2X1M U349 (.Y(n289), 
	.B1(n158), 
	.B0(n358), 
	.A1N(n158), 
	.A0N(\memory[12][6] ));
   OAI2BB2X1M U350 (.Y(n290), 
	.B1(n158), 
	.B0(n357), 
	.A1N(n158), 
	.A0N(\memory[12][7] ));
   OAI2BB2X1M U351 (.Y(n291), 
	.B1(n160), 
	.B0(n364), 
	.A1N(n160), 
	.A0N(\memory[13][0] ));
   OAI2BB2X1M U352 (.Y(n292), 
	.B1(n160), 
	.B0(n363), 
	.A1N(n160), 
	.A0N(\memory[13][1] ));
   OAI2BB2X1M U353 (.Y(n293), 
	.B1(n160), 
	.B0(n362), 
	.A1N(n160), 
	.A0N(\memory[13][2] ));
   OAI2BB2X1M U354 (.Y(n294), 
	.B1(n160), 
	.B0(n361), 
	.A1N(n160), 
	.A0N(\memory[13][3] ));
   OAI2BB2X1M U355 (.Y(n295), 
	.B1(n160), 
	.B0(n360), 
	.A1N(n160), 
	.A0N(\memory[13][4] ));
   OAI2BB2X1M U356 (.Y(n296), 
	.B1(n160), 
	.B0(n359), 
	.A1N(n160), 
	.A0N(\memory[13][5] ));
   OAI2BB2X1M U357 (.Y(n297), 
	.B1(n160), 
	.B0(n358), 
	.A1N(n160), 
	.A0N(\memory[13][6] ));
   OAI2BB2X1M U358 (.Y(n298), 
	.B1(n160), 
	.B0(n357), 
	.A1N(n160), 
	.A0N(\memory[13][7] ));
   OAI2BB2X1M U359 (.Y(n299), 
	.B1(n161), 
	.B0(n364), 
	.A1N(n161), 
	.A0N(\memory[14][0] ));
   OAI2BB2X1M U360 (.Y(n300), 
	.B1(n161), 
	.B0(n363), 
	.A1N(n161), 
	.A0N(\memory[14][1] ));
   OAI2BB2X1M U361 (.Y(n301), 
	.B1(n161), 
	.B0(n362), 
	.A1N(n161), 
	.A0N(\memory[14][2] ));
   OAI2BB2X1M U362 (.Y(n302), 
	.B1(n161), 
	.B0(n361), 
	.A1N(n161), 
	.A0N(\memory[14][3] ));
   OAI2BB2X1M U363 (.Y(n303), 
	.B1(n161), 
	.B0(n360), 
	.A1N(n161), 
	.A0N(\memory[14][4] ));
   OAI2BB2X1M U364 (.Y(n304), 
	.B1(n161), 
	.B0(n359), 
	.A1N(n161), 
	.A0N(\memory[14][5] ));
   OAI2BB2X1M U365 (.Y(n305), 
	.B1(n161), 
	.B0(n358), 
	.A1N(n161), 
	.A0N(\memory[14][6] ));
   OAI2BB2X1M U366 (.Y(n306), 
	.B1(n161), 
	.B0(n357), 
	.A1N(n161), 
	.A0N(\memory[14][7] ));
   OAI2BB2X1M U367 (.Y(n307), 
	.B1(n163), 
	.B0(n364), 
	.A1N(n163), 
	.A0N(\memory[15][0] ));
   OAI2BB2X1M U368 (.Y(n308), 
	.B1(n163), 
	.B0(n363), 
	.A1N(n163), 
	.A0N(\memory[15][1] ));
   OAI2BB2X1M U369 (.Y(n309), 
	.B1(n163), 
	.B0(n362), 
	.A1N(n163), 
	.A0N(\memory[15][2] ));
   OAI2BB2X1M U370 (.Y(n310), 
	.B1(n163), 
	.B0(n361), 
	.A1N(n163), 
	.A0N(\memory[15][3] ));
   OAI2BB2X1M U371 (.Y(n311), 
	.B1(n163), 
	.B0(n360), 
	.A1N(n163), 
	.A0N(\memory[15][4] ));
   OAI2BB2X1M U372 (.Y(n312), 
	.B1(n163), 
	.B0(n359), 
	.A1N(n163), 
	.A0N(\memory[15][5] ));
   OAI2BB2X1M U373 (.Y(n313), 
	.B1(n163), 
	.B0(n358), 
	.A1N(n163), 
	.A0N(\memory[15][6] ));
   OAI2BB2X1M U374 (.Y(n314), 
	.B1(n163), 
	.B0(n357), 
	.A1N(n163), 
	.A0N(\memory[15][7] ));
   INVX2M U375 (.Y(n341), 
	.A(N12));
   AO21XLM U376 (.Y(n186), 
	.B0(n365), 
	.A1(n166), 
	.A0(RdData_VLD));
   DLY1X4M U377 (.Y(n370), 
	.A(test_se));
   DLY1X4M U378 (.Y(n371), 
	.A(test_se));
   DLY1X4M U379 (.Y(n372), 
	.A(test_se));
   DLY1X4M U380 (.Y(n373), 
	.A(test_se));
endmodule


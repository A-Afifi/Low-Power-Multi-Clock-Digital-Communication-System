// ************************************************************* //
//                      Module : Integer_ClkDiv_tb               //
//                      Author : Ahmed_Afifi                     //
// ************************************************************* //

`timescale 1ns/1ps

module Integer_ClkDiv_tb ();

//******************************* Parameters *******************************
parameter   ratio_Width_tb = 8 ,
            ref_clk_PERIOD = 2 ;  // 500 MHz

//******************************* DUT Signals ******************************

reg                             i_ref_clk_tb;
reg                             i_rst_n_tb;
reg                             i_clk_en_tb;
reg    [ratio_Width_tb-1:0]     i_dev_ratio_tb;
wire                            o_div_clk_tb;

//***************************** DUT Instantation ****************************
Integer_ClkDiv #(.ratio_Width(ratio_Width_tb)) DUT (
.i_ref_clk(i_ref_clk_tb),
.i_rst_n(i_rst_n_tb),
.i_clk_en(i_clk_en_tb),
.i_dev_ratio(i_dev_ratio_tb),
.o_div_clk(o_div_clk_tb)
);


//******************************* initial block *******************************
initial 
begin
    // System Functions
    $dumpfile("Int_ClkDiv_DUMP.vcd") ;       
    $dumpvars; 

    // initialization
    initialize() ;
    // Reset 
    #10;
    reset();

    //////////////////////////////////////////////////////////////// Name Print /////////////////////////////////////////////////////////////////////
    $display("\nName : Ahmed Mohamed Afifi");
    $display("Name : Integer_ClkDiv\n\n");


    #10;
    @(posedge i_ref_clk_tb);
    //////////////////////////////////////////////////////////////// Test Case (1) /////////////////////////////////////////////////////////////////////
    Test_Case_num('d1);
    $display("Dividing by 8 \n");
    Freq_Div_Op('d8);


    #10;
    @(posedge i_ref_clk_tb);
    //////////////////////////////////////////////////////////////// Test Case (2) /////////////////////////////////////////////////////////////////////
    Test_Case_num('d2);
    $display("Dividing by 5 \n");
    Freq_Div_Op('d5);
    

    #10;
    @(posedge i_ref_clk_tb) ;
    //////////////////////////////////////////////////////////////// Test Case (3) /////////////////////////////////////////////////////////////////////
    Test_Case_num('d3);
    $display("Dividing by 1 \n");
    Freq_Div_Op('d1);


    #10;
    @(posedge i_ref_clk_tb) ;
    //////////////////////////////////////////////////////////////// Test Case (4) /////////////////////////////////////////////////////////////////////
    Test_Case_num('d4);
    $display("Dividing by 0 \n");
    Freq_Div_Op('d0);


    #10;
    @(posedge i_ref_clk_tb) ;
    //////////////////////////////////////////////////////////////// Test Case (5) /////////////////////////////////////////////////////////////////////
    Test_Case_num('d5);
    $display("Dividing by 127 \n");
    Freq_Div_Op('d127);


    #10;
    @(posedge i_ref_clk_tb) ;
    //////////////////////////////////////////////////////////////// Test Case (6) /////////////////////////////////////////////////////////////////////
    Test_Case_num('d6);
    $display("Dividing by 255 \n");
    Freq_Div_Op('d255);


    #10;
    @(posedge i_ref_clk_tb) ;
    //////////////////////////////////////////////////////////////// Test Case (7) /////////////////////////////////////////////////////////////////////
    Test_Case_num('d7);
    $display("From high i_dev_ratio to low corner case \n");

    i_dev_ratio_tb       =  'd8 ;
    i_clk_en_tb          = 1'b1;   

    repeat (8) @(posedge i_ref_clk_tb);
    repeat (10) @(posedge i_ref_clk_tb); 
    @(negedge i_ref_clk_tb); 
    
    i_dev_ratio_tb       =  'd4 ;

    repeat (15) @(posedge i_ref_clk_tb); 
    #20 ;
    i_clk_en_tb          = 1'b0; 



    
    #100;
    $stop ;

end    

 

//*************************************************************************************************************************************************//
//***************************************************************** TASKS *************************************************************************//
//*************************************************************************************************************************************************//


//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//******************************************************** Test_Case_num *******************************************//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
task Test_Case_num ;
    input [5:0] num ;
  begin
        $write ("Test Case (%d ) : ",num);
  end
endtask



//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//**************************************************** Signals Initialization **************************************//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
task initialize ;
  begin
	i_ref_clk_tb         = 1'b0;
	i_rst_n_tb           = 1'b1;    
	i_clk_en_tb          = 1'b0;   
	i_dev_ratio_tb       =  'd4;

  end
endtask


//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//************************************************* RESET **********************************************************//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
task reset ;
    begin
        i_rst_n_tb  = 1'b1;
        @(posedge i_ref_clk_tb);
        i_rst_n_tb  = 1'b0;
        #40;
        @(negedge i_ref_clk_tb);
        i_rst_n_tb  = 1'b1;
    end
endtask

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//************************************************* Freq_Div_Op ****************************************************//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
task Freq_Div_Op ;
    input [ratio_Width_tb-1:0] div_ratio ;
    begin 
        i_dev_ratio_tb       =  div_ratio ;
        i_clk_en_tb          = 1'b1;   
        #510 ;
        @(posedge i_ref_clk_tb); 
        i_clk_en_tb          = 1'b0; 
        @(posedge i_ref_clk_tb); 
    end
endtask


//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//******************************************************* Clock Generator ******************************************//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
always #(ref_clk_PERIOD/2) i_ref_clk_tb = ~i_ref_clk_tb ;



endmodule
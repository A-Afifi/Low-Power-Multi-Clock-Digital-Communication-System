

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO SYS_TOP 
  PIN SI[3] 
    ANTENNAPARTIALMETALAREA 1.827 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.78787 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 6.641 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.1356 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 7.885 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.1193 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 237.348 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1151.82 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA45 ;
  END SI[3]
  PIN SI[2] 
    ANTENNAPARTIALMETALAREA 6.054 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.1197 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 29.624 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 142.684 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 12.135 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 58.5618 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 292.189 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1419.21 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END SI[2]
  PIN SI[1] 
    ANTENNAPARTIALMETALAREA 4.605 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.1501 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 19.588 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 94.4107 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.131 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 39.3025 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 193.164 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 939.298 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 3.38649 LAYER VIA45 ;
  END SI[1]
  PIN SI[0] 
    ANTENNAPARTIALMETALAREA 0.405 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.94805 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 9.689 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.7965 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 208.83 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 1011.04 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA34 ;
  END SI[0]
  PIN SO[3] 
    ANTENNADIFFAREA 0.537 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.611 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.74891 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 54.5245 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 260.697 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.53405 LAYER VIA34 ;
  END SO[3]
  PIN SO[2] 
    ANTENNADIFFAREA 0.537 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 23.101 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 111.308 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1274 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 186.836 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 898.785 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.850078 LAYER VIA34 ;
  END SO[2]
  PIN SO[1] 
    ANTENNAPARTIALMETALAREA 4.273 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.5531 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.168 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.00048 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 32.002 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 154.122 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 181.66 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 874.832 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.0241 LAYER VIA56 ;
  END SO[1]
  PIN SO[0] 
    ANTENNAPARTIALMETALAREA 2.85 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.7085 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 200.693 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 966.54 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.07233 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.268 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48148 LAYER METAL4 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 203.77 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 983.549 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.90126 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 44.188 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 212.737 LAYER METAL5 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 711.095 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 3425.99 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.90126 LAYER VIA56 ;
  END SO[0]
  PIN scan_clk 
    ANTENNAPARTIALMETALAREA 0.255 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.22655 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.81 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.632 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.23232 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 0.574507 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 2.90913 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END scan_clk
  PIN scan_rst 
    ANTENNAPARTIALMETALAREA 1.517 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.29677 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 13.739 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.277 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.2166 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 22.934 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 110.89 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1599 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 258.887 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1252.61 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 3.38649 LAYER VIA45 ;
  END scan_rst
  PIN test_mode 
    ANTENNAPARTIALMETALAREA 2.665 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.8187 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 32.0482 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 153.148 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.414466 LAYER VIA23 ;
  END test_mode
  PIN SE 
    ANTENNAPARTIALMETALAREA 1.421 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.83501 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1755 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 8.9265 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 42.1607 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.205698 LAYER VIA23 ;
  END SE
  PIN RST_N 
    ANTENNAPARTIALMETALAREA 0.729 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.50649 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.268 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48148 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 12.641 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 60.9956 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 321.52 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1553.87 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 3.38649 LAYER VIA45 ;
  END RST_N
  PIN UART_CLK 
    ANTENNAPARTIALMETALAREA 0.241 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.15921 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.862 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.14862 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.412 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.9865 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 0.969897 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 4.87377 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END UART_CLK
  PIN REF_CLK 
    ANTENNAPARTIALMETALAREA 0.537 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.58297 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.076 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.798 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 1.46585 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 7.13366 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END REF_CLK
  PIN UART_RX_IN 
    ANTENNAPARTIALMETALAREA 0.669 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.21789 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 8.28 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.2116 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2483 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 57.025 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 275.112 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.65786 LAYER VIA34 ;
  END UART_RX_IN
  PIN UART_TX_O 
    ANTENNADIFFAREA 0.524 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.975 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3098 LAYER METAL3 ;
  END UART_TX_O
  PIN parity_error 
    ANTENNAPARTIALMETALAREA 29.27 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 140.789 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.124 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.59884 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 19.046 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 91.8037 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 509.037 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2462.25 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 4.06379 LAYER VIA56 ;
  END parity_error
  PIN framing_error 
    ANTENNAPARTIALMETALAREA 44.13 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 212.265 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNADIFFAREA 0.6 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 5.238 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 25.3872 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 112.639 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 551.971 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END framing_error
END SYS_TOP

END LIBRARY
